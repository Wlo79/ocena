��-     �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�	estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.2.2�ub�n_estimators�K(�estimator_params�(hhhhhhhhhht��base_estimator��
deprecated��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        hKhNhG        hG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK*��h*�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�class_number��learning_time��learning_intensity��from_coursebook��from_notebook��from_many_notebooks��	from_apps��from_websites��from_flashards��
from_books��prosGoodMark��prosInterest��prosPositivMark��prosJoy��prosJob��prosStudies��prosNone��badWellBeing��busySchedule��hatred_to_subject��entertainment��richSocialLife��badFactorsNone��goodAttitude��determination��goodSchedule��goodScheduleLearn��joyResignation��goodFactorsNone��actual_motivation��gradePredictions��subject_grad��subject_other��subject_prof��teacher_behaviour_inert��teacher_behaviour_normal��teacher_behaviour_watch��questions_notSurprised��questions_surprised��sex_man��sex_notGiven��	sex_woman�et�b�n_features_in_�K*�
n_outputs_�K�classes_�h)h,K ��h.��R�(KK��h3�i8�����R�(K�<�NNNJ����J����K t�b�C0                                          �t�b�
n_classes_�K�
estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hKhNhJ�
hG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h3�f8�����R�(KhoNNNJ����J����K t�b�C0              �?       @      @      @      @�t�bhsh'�scalar���hnC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hK�
node_count�K��nodes�h)h,K ��h.��R�(KK���h3�V56�����R�(Kh7N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(h�hnK ��h�hnK��h�hnK��h�hK��h�hK ��h�hnK(��h�hK0��uK8KKt�b�B�$         f       &             �?�<U����?�            `u@       5                    @v�f��?y            `g@                           �?�wvJ;�??            �V@                           @pƵHPS�?             :@       
                    �?     ��?             0@                           �?@4և���?	             ,@������������������������       �                     (@       	                    �?      �?              @������������������������       �                     �?������������������������       �                     �?                           �?      �?              @������������������������       �                     �?������������������������       �                     �?                           �?H�z�G�?             $@                           �?      �?              @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @       *       
             �?     d�?-             P@                           �?v���n(�?            �@@                           �?P���� �?             7@                           @�lO���?             3@                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     0@                           �?      �?             @������������������������       �                      @������������������������       �                      @        #                    �?p=
ףp�?             $@!       "                    �?      �?             @������������������������       �                     @������������������������       �                     �?$       )       )             �?�q�q�?             @%       &                    �?      �?             @������������������������       �                     �?'       (                     �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @+       0                    �?��b�=�?             ?@,       /                    @      �?             8@-       .       )             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     6@1       2                    �?:/����?             @������������������������       �                      @3       4       '             �?���Q��?             @������������������������       �                      @������������������������       �                     @6       _                    �?x��;���?:            @X@7       Z                    �?Vw�����?3            @U@8       K                    �?�������?/            �S@9       F                    @|� \4(�?            �B@:       C                    @��t��L�?             ?@;       B                    @�GN�z�?             6@<       A                    �?�eP*L��?             &@=       @       '             �?�q�q�?             "@>       ?                     �?      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     &@D       E       )             �?X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @G       H                    �?�q�q�?             @������������������������       �                     �?I       J                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?L       M                    �?�p ��?            �D@������������������������       �                     @N       U       	             �?b�h�d.�?            �A@O       T       "             �?�>����?             ;@P       Q                    �? ��WV�?             :@������������������������       �                     5@R       S                    @z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?V       W                    �?      �?              @������������������������       �                      @X       Y                    �?�q�q�?             @������������������������       �                     @������������������������       �                      @[       \                    @:/����?             @������������������������       �                     @]       ^       #             �?      �?             @������������������������       �                      @������������������������       �                      @`       c                    @      �?             (@a       b                    @r�q��?             @������������������������       �                     @������������������������       �                     �?d       e                    �?�q�q�?             @������������������������       �                      @������������������������       �                     @g       �                    �?�c�Ę�?_            `c@h       k                    �?���#���?9             V@i       j                    �?      �?
             0@������������������������       �        	             .@������������������������       �                     �?l       q                     �?�%���^�?/             R@m       p                    �?8�Z$���?             *@n       o                    �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @r       �                    �?��;F���?(            �M@s       �                    �?�q-74��?%            �K@t       u                    �?`՟�G��?             ?@������������������������       �        	             (@v       �       $             �?�d�����?             3@w       �                    �?�q�q�?	             (@x       �       !             �?���|���?             &@y       �                    @�<ݚ�?             "@z              )             �?      �?              @{       ~       "             �?r�q��?             @|       }                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �? �q�q�?             8@�       �                    �?r�q��?             @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     2@�       �       
             �?      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �?����cZ�?&            �P@�       �                    �?�q�q�?             ;@�       �                    �?      �?             4@������������������������       �                     @�       �                    @      �?
             0@������������������������       �                     (@�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @�       �       #             �?և���X�?             @������������������������       �                      @�       �                    �?z�G�z�?             @������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �       !             �?�G�z��?             D@�       �                    �?�	j*D�?             :@������������������������       �                     &@�       �                    @��S���?	             .@�       �                    �?�<ݚ�?             "@�       �                    �?      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     ,@�t�b�values�h)h,K ��h.��R�(KK�KK��h�B�        F@     �J@     �R@     @U@     �O@      6@      @      @      ?@      N@     �O@      6@      @      @      ?@     �G@      �?                       @      0@      @      �?                       @      *@      �?                              �?      *@                                              (@                                      �?      �?                                              �?                                      �?                                              �?              �?                              �?                                                              �?                                      @      @      �?                              �?      @      �?                              �?              �?                              �?                                                              �?                                      @                                       @                              @      @      .@      D@                      @      �?      &@      0@                      @              @      0@                      �?               @      0@                      �?               @                                               @                              �?                                                                      0@                       @               @                                               @                               @                                               @      �?      @                                      �?      @                                              @                                      �?                                       @              @                               @               @                                              �?                               @              �?                                              �?                               @                                                               @                              �?       @      @      8@                      �?              �?      6@                      �?              �?                              �?                                                              �?                                                      6@                               @      @       @                               @                                                      @       @                                               @                                      @                                                      *@      O@      6@                               @      N@      1@                              @      M@      .@                              @      7@      "@                              @      5@      @                              @      1@                                      @      @                                      @      @                                      @      @                                      @                                                      @                                              @                                       @                                                      &@                                              @      @                                      @                                                      @                                       @      @                                      �?                                              �?      @                                              @                                      �?                                             �A@      @                                      @                                              =@      @                                      9@       @                                      9@      �?                                      5@                                              @      �?                                      @                                                      �?                                              �?                                      @      @                                               @                                      @       @                                      @                                                       @                              @       @       @                              @                                                       @       @                                               @                                       @                                      @       @      @                              @              �?                              @                                                              �?                                       @      @                                       @                                                      @      C@      H@      F@      9@                      =@      >@      :@      @                      .@      �?                                      .@                                                      �?                                      ,@      =@      :@      @                              &@       @                                      @       @                                      @                                                       @                                       @                                      ,@      2@      8@      @                      ,@      2@      7@                              ,@      1@                                              (@                                      ,@      @                                      @      @                                      @      @                                      @       @                                      @      �?                                      @      �?                                       @      �?                                              �?                                       @                                              @                                               @                                                      �?                                               @                                              �?                                      @                                                      �?      7@                                      �?      @                                      �?       @                                      �?                                                       @                                              @                                              2@                                              �?      @                                      �?                                                      @                      "@      2@      2@      6@                      "@      2@                                      @      .@                                      @                                              �?      .@                                              (@                                      �?      @                                      �?                                                      @                                      @      @                                               @                                      @      �?                                      @                                              �?      �?                                      �?                                                      �?                                                      2@      6@                                      2@       @                                      &@                                              @       @                                      @       @                                      @      �?                                      @                                                      �?                                              �?                                              @                                              ,@                �t�bubhhubh)��}�(hhhhhNhKhKhG        hKhNhJ/��hG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKׅ�h��B/         �                    @���;R��?�            `u@       e       
             �?�L��P��?�            `o@       <                    �?(�T����?f             c@                           �?������?=            �V@                           �?�e����?            �C@������������������������       �        
             *@                           �?ȵHPS!�?             :@       	                    �?�X�<ݺ?             2@������������������������       �                     "@
                           �?�����H�?             "@������������������������       �                     @                            @�q�q�?             @������������������������       �                     �?                           @      �?              @������������������������       �                     �?������������������������       �                     �?              #             �?      �?              @                           @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @       7       )             �?��m���?!             J@       6                    �?     ��?             @@       '       &             �?<+	���?             >@                            @4և����?	             ,@              #             �?      �?             @������������������������       �                      @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?       $       "             �?ffffff�?             $@        !                    �?z�G�z�?             @������������������������       �                     �?"       #                    �?      �?             @������������������������       �                     @������������������������       �                     �?%       &                    �?���Q��?             @������������������������       �                      @������������������������       �                     @(       -                    �?     ��?             0@)       *                    �?��!pc�?             &@������������������������       �                     �?+       ,                    @ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?.       5                    �?���Q��?             @/       0                    �?      �?             @������������������������       �                     �?1       4                    @�q�q�?             @2       3                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @8       ;       #             �?ףp=
�?
             4@9       :                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     1@=       X                     @]"?ӧ
�?)             O@>       Q                    �?�ѷQC�?            �B@?       J                    �?V}��b�?             9@@       C                    �?�eP*L��?	             &@A       B       )             �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?D       I       )             �?�q�q�?             @E       H                    �?�q�q�?             @F       G                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @K       L                    @N��)x9�?
             ,@������������������������       �                     @M       N                    @X�<ݚ�?             "@������������������������       �                     @O       P       &             �?r�q��?             @������������������������       �                     @������������������������       �                     �?R       W                    �?r�q��?             (@S       T                     �?�8��8��?             @������������������������       �                     @U       V       #             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @Y       `                    @b2U0*��?             9@Z       _                     �?      �?              @[       \                    �?؇���X�?             @������������������������       �                     @]       ^                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?a       d                    �?������?
             1@b       c                    �?@4և���?             ,@������������������������       �                     *@������������������������       �                     �?������������������������       �                     @f       �                    �?2M���c�?<            �X@g       �       "             �?��8�l�?"            �J@h       �       &             �?l]?���?            �F@i       x                    �?�q-��?             :@j       k                    �?H�7�&��?	             .@������������������������       �                     �?l       u                    �?����S�?             ,@m       t                    �?�C��2(�?             &@n       s                    �?؇���X�?             @o       p                    @z�G�z�?             @������������������������       �                      @q       r                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @v       w       $             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @y       �                    �?���!pc�?             &@z       }                    @B{	�%��?             "@{       |                    �?���Q��?             @������������������������       �                      @������������������������       �                     @~                           @      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @�       �                    �?���y4F�?             3@�       �                    @�t����?	             1@�       �       )             �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     *@������������������������       �                      @�       �                    �?      �?              @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?����?�?            �F@�       �       $             �?      �?              @������������������������       �                     @�       �                     �?���Q��?             @������������������������       �                      @������������������������       �                     @�       �                    �?��o^_�?            �B@�       �                    �?&%�ݒ��?             5@�       �                    @և���X�?             @�       �                    �?z�G�z�?             @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                      @�       �       $             �?@4և���?             ,@������������������������       �                     *@������������������������       �                     �?�       �       "             �?     @�?	             0@�       �                     @x9/���?             ,@������������������������       �                     @�       �                    �?      �?              @������������������������       �                     @�       �                    �?�Q����?             @�       �                    �?      �?             @�       �                     @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �       %             �?ą�l��?6            �V@�       �                    �?|�ʒ���?             3@������������������������       �                     (@�       �                    @����>4�?             @�       �       '             �?      �?             @������������������������       �                      @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �       !             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    @�[��"e�?*             R@�       �                    @��X��?#             L@�       �                     @r�q��?
             (@������������������������       �                     �?�       �                    �?"pc�
�?	             &@������������������������       �                     @�       �                    �?      �?             @������������������������       �                     �?�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?�GN�z�?             F@�       �                    �?���N8�?             5@������������������������       �                     4@������������������������       �                     �?�       �                    @�û��|�?             7@�       �                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    �?������?
             1@�       �       	             �?     ��?	             0@�       �                    @�r����?             .@������������������������       �                     *@������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                    @     ��?             0@������������������������       �                     @������������������������       �                     &@�t�bh�h)h,K ��h.��R�(KK�KK��h�BP(        ;@     �H@     @W@      S@      P@     �@@      :@      H@     �V@      K@      7@      $@      7@     �B@     �J@      8@      $@      @      0@      :@     �@@      @      @      @      0@      7@                                      *@                                              @      7@                                      �?      1@                                              "@                                      �?       @                                              @                                      �?       @                                              �?                                      �?      �?                                      �?                                                      �?                                       @      @                                       @      �?                                              �?                                       @                                                      @                                              @     �@@      @      @      @              @      .@      @      @      @              @      .@      @      @      @              �?      @      @      @      @              �?       @      �?                                       @                                      �?              �?                              �?                                                              �?                                      �?       @      @      @                      �?              @                                              �?                              �?              @                                              @                              �?                                                       @              @                               @                                                              @               @      (@              �?      �?                      "@              �?      �?                                              �?                      "@              �?                              "@                                                              �?                       @      @                                       @       @                                      �?                                              �?       @                                      �?      �?                                      �?                                                      �?                                              �?                                              �?                                                       @                                      2@                       @                      �?                       @                                               @                      �?                                              1@                              @      &@      4@      3@      @              @      @      ,@      @      @              @      @      @      @      @              @      @                                      @      �?                                      @                                                      �?                                       @      @                                       @      �?                                      �?      �?                                      �?                                                      �?                                      �?                                                      @                                                      @      @      @                              @                                                      @      @                                      @                                              �?      @                                              @                                      �?                      �?              "@       @                      �?              @       @                                      @                              �?                       @                                               @                      �?                                                              @                                      @      @      *@                              @       @                                      @      �?                                      @                                              �?      �?                                              �?                                      �?                                                      �?                                              @      *@                                      �?      *@                                              *@                                      �?                                              @                              @      &@     �B@      >@      *@      @              @      >@       @      @      @              @      =@      @      @       @               @      ,@      @      @       @                      (@      �?       @                                              �?                              (@      �?      �?                              $@      �?                                      @      �?                                      @      �?                                       @                                               @      �?                                              �?                                       @                                               @                                              @                                               @              �?                                              �?                               @                                       @       @      @       @       @               @              @       @       @               @              @                               @                                                              @                                                       @       @                                       @                                                       @                       @                                      @      .@                                       @      .@                                       @       @                                       @                                                       @                                              *@                                       @                                                      �?      @       @      �?                              @       @                                               @                                      @                                      �?                      �?                                              �?                      �?                              @      @      @      6@      @      �?      @      @                                              @                                      @       @                                               @                                      @                                                              @      6@      @      �?                      @      1@      �?                              @      @                                      �?      @                                      �?       @                                      �?                                                       @                                               @                                       @                                                      *@      �?                                      *@                                                      �?                              @      @      @      �?                      @      @      @      �?                                      @                              @      @              �?                      @                                              �?      @              �?                      �?      @                                      �?      �?                                              �?                                      �?                                                       @                                                              �?                               @                      �?      �?      @      6@     �D@      7@              �?      @      *@               @                              (@                              �?      @      �?               @              �?      @                                               @                                      �?      �?                                              �?                                      �?                                                              �?               @                              �?                                                               @      �?                      "@     �D@      5@      �?                      "@      B@      $@      �?                      "@       @              �?                                                                      "@       @                                      @                                               @       @                                      �?                                              �?       @                                      �?                                                       @                                              A@      $@                                      4@      �?                                      4@                                                      �?                                      ,@      "@                                      �?      @                                              @                                      �?                                              *@      @                                      *@      @                                      *@       @                                      *@                                                       @                                              �?                                              �?                                      @      &@                                      @                                                      &@�t�bubhhubh)��}�(hhhhhNhKhKhG        hKhNhJu�7hG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK˅�h��Bh,         \       %             �?�G-,�?�            `u@       %                     @�G�z��?b            �b@                           �?߼�xV4�?)             N@                           �?�lg����?            �E@������������������������       �                     @                           �?�G�z�?             D@                           �?�	j*D�?            �C@                           �?     ��?             @@	                           @���|���?	             &@
                           �?�<ݚ�?             "@������������������������       �                     �?                           �?      �?              @������������������������       �                     @                            @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @                            �?�����?             5@                           �?8�Z$���?             *@������������������������       �                     $@                           �?�q�q�?             @������������������������       �                     �?              !             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @              #             �?؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?       $                    �?f�t���?             1@        #                    �?p=
ףp�?             $@!       "                    �?      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @&       )                    �?��� Ce�?9            �V@'       (                    �?     ��?             0@������������������������       �                     *@������������������������       �                     @*       7                    �?�6<�v$�?1            �R@+       6                    @H�z�G�?             4@,       1       #             �?H�7�&��?             .@-       0                    �?VUUUUU�?             @.       /                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?2       5                    �?�8��8��?	             (@3       4                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     "@������������������������       �                     @8       [                    �?�
��?              K@9       X                    �?~e�.y0�?             J@:       O                    �?6�G�ܸ�?             G@;       D                    @x�W��#�?             7@<       C                    @B{	�%��?             "@=       B                    �?      �?              @>       A                     @؇���X�?             @?       @                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     �?E       N                    �?      �?             ,@F       M                    �?�q�q�?             (@G       L       "             �?����X�?             @H       K                    �?���Q��?             @I       J       $             �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @P       S                    �?$G�h��?             7@Q       R                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?T       U                    �?P���Q�?             4@������������������������       �                     ,@V       W                    �?r�q��?             @������������������������       �                     �?������������������������       �                     @Y       Z       '             �?r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @]       �                    @�8��8��?q             h@^       �       
             �?�j;��W�?;            �V@_       ~                    �?L䯦s#�?!            �J@`       s                    @,W�k^�?            �D@a       h                    �?�l'l��?             ?@b       g                    �?      �?              @c       d                    �?z�G�z�?             @������������������������       �                      @e       f                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @i       r                    �?8����?             7@j       q                    �?��
ц��?             *@k       p                    �?�z�G��?             $@l       o                    �?      �?             @m       n                    @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     $@t       }                    �?ffffff�?             $@u       x                     �?      �?              @v       w                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @y       z                     �?VUUUUU�?             @������������������������       �                     �?{       |                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @       �                    �?�������?	             (@������������������������       �                     �?�       �                    �?�C��2(�?             &@������������������������       �                     @�       �                    @r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                    �?��I!��?            �B@�       �                    �?ȵHPS!�?             :@�       �                    @P���Q�?             4@������������������������       �        	             *@�       �                    �?؇���X�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �       #             �?�q�q�?             @������������������������       �                      @�       �                     �?      �?             @������������������������       �                      @������������������������       �                      @�       �                    �?��!pc�?             &@�       �                    �?      �?              @�       �                    �?z�G�z�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �?j���� �?6            �Y@�       �                    �?�F_��C�?             M@�       �                    @�{���w�?            �F@�       �                    @���	7I�?            �C@�       �       (             �?��J���?             6@�       �                     �?&%�ݒ��?
             5@�       �                    �?      �?             (@������������������������       �                     �?�       �                    @"pc�
�?             &@�       �       
             �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �       
             �?�����H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     1@�       �       #             �?�8��8��?             @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �?��WV��?             *@�       �                    �?{�G�z�?             $@�       �       #             �?z�G�z�?             @������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                    @�eP*L��?             F@������������������������       �                     5@�       �       )             �?�LQ�1	�?             7@�       �                    �?�θ�?             *@�       �                    �?      �?              @�       �                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     $@�t�bh�h)h,K ��h.��R�(KK�KK��h�B&        D@     �L@      N@     @T@     @R@      ?@      A@     �J@      D@      0@       @      @      0@      ;@      @       @       @              0@      ;@                                      @                                              *@      ;@                                      (@      ;@                                      @      :@                                      @      @                                       @      @                                      �?                                              �?      @                                              @                                      �?       @                                      �?                                                       @                                       @                                               @      3@                                       @      &@                                              $@                                       @      �?                                      �?                                              �?      �?                                              �?                                      �?                                                       @                                      @      �?                                      @                                                      �?                                      �?                                                              @       @       @                              @      �?       @                              @      �?                                      @                                                      �?                                                       @                                      @                      2@      :@     �@@       @              @      *@                                      @      *@                                                                                      @      @      :@     �@@       @               @       @      (@      @                               @      (@      �?                              �?      �?      �?                              �?      �?                                      �?                                                      �?                                                      �?                              �?      &@                                      �?       @                                      �?                                                       @                                              "@                                                      @                              @      ,@      ;@       @               @      @      ,@      ;@       @                       @      "@      ;@       @                      �?      @       @      @                      �?      @      �?                              �?      @                                      �?      @                                      �?      �?                                      �?                                                      �?                                              @                                              �?                                                      �?                                              @      @                                      @      @                                       @      @                                       @      @                                      �?      @                                              @                                      �?                                              �?                                                       @                                      @                                                       @                      �?       @      3@      �?                      �?       @                                               @                                      �?                                                              3@      �?                                      ,@                                              @      �?                                              �?                                      @                              �?      @                                      �?                                                      @                                                                               @      @      @      4@     @P@     �Q@      :@      @      @      4@     �L@      @              @      @      0@      =@                      @      @      .@      3@                              �?      ,@      0@                              �?      @                                      �?      @                                               @                                      �?       @                                               @                                      �?                                                      @                                              @      0@                                      @      @                                      @      @                                      @      @                                      @      �?                                      @                                                      �?                                               @                                      @                                                      @                                              $@                      @       @      �?      @                      @       @      �?      �?                      @      �?                                              �?                                      @                                                      �?      �?      �?                                      �?                                      �?              �?                                              �?                              �?                                                               @                              �?      �?      $@                              �?                                                      �?      $@                                              @                                      �?      @                                      �?                                                      @                       @              @      <@      @                                      7@      @                                      3@      �?                                      *@                                              @      �?                                      �?      �?                                              �?                                      �?                                              @                                              @       @                                       @                                               @       @                                       @                                                       @               @              @      @                       @              �?      @                                      �?      @                                      �?      �?                                      �?                                                      �?                                              @                       @                      �?                       @                                                                      �?                                      @                                                       @      Q@      :@                               @      F@      @                              @     �B@       @                              @      A@      �?                              @      1@      �?                              @      1@      �?                              @      "@                                      �?                                               @      "@                                       @      @                                              @                                       @                                                      @                                               @      �?                                              �?                                       @                                      �?                                                      1@                                       @      @      �?                               @              �?                                              �?                               @                                                      @                                       @      @      @                               @      @      @                                      @      �?                                      @                                              �?      �?                                              �?                                      �?                                       @              @                               @                                                              @                                      @                                              8@      4@                                      5@                                              @      4@                                      @      $@                                      @      @                                      �?      @                                              @                                      �?                                               @                                                      @                                              $@�t�bubhhubh)��}�(hhhhhNhKhKhG        hKhNhJ��!XhG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKㅔh��B�1         �                    @��k��?�            `u@       A                    �?*��Ӥ��?�             h@       ,                    �?��Ϭ&�?K            �[@                           @���W�?/            �Q@       
                    �?K&:~��?             3@              '             �?ףp=
�?             $@������������������������       �                      @       	                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@              
             �?R�k���?!            �I@                           @�q�q�?             8@                           �?�����?             5@                           �?      �?              @������������������������       �                     �?������������������������       �                     �?                           �?�}�+r��?             3@������������������������       �                     ,@                           �?z�G�z�?             @              "             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @       %                    @���'���?             ;@                             �?     ��?             0@                             @8�Z$���?             *@������������������������       �                     @                           �?�<ݚ�?             "@������������������������       �                     @������������������������       �                      @!       $                    �?VUUUUU�?             @"       #                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?&       +                    @�eP*L��?             &@'       *                    �?X�<ݚ�?             "@(       )                    �?r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @-       2                    �?>
ףp=�?             D@.       1                    �?X�<ݚ�?             "@/       0       %             �?����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @3       @                    @��b�=�?             ?@4       5                    �?
�b�m��?             =@������������������������       �                     .@6       7       %             �?      �?	             ,@������������������������       �                     @8       ?       (             �?���(\��?             $@9       >                     @�$I�$I�?             @:       =                    �?�q�q�?             @;       <                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @B       g                    �?� t���?6            �T@C       Z                    �?!�$|�*�?            �F@D       K                    �?     ��?             @@E       F       #             �?      �?              @������������������������       �                     @G       J                    �?�q�q�?             @H       I                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?L       U       $             �?��8��8�?             8@M       P                    �?ffffff�?             4@N       O                    @�IєX�?             1@������������������������       �                     0@������������������������       �                     �?Q       T       )             �?VUUUUU�?             @R       S                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?V       W                    �?      �?             @������������������������       �                      @X       Y                    �?      �?              @������������������������       �                     �?������������������������       �                     �?[       b                    �?����W�?	             *@\       a                    �?{�G�z�?             @]       `       #             �?      �?             @^       _       %             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?c       f       '             �?      �?              @d       e                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @h       w                    @u#����?             C@i       j                    �?П[;U��?             =@������������������������       �        	             0@k       t                    �?޾�z�<�?             *@l       m       #             �?z�G�z�?             $@������������������������       �                     �?n       o                     @�����H�?             "@������������������������       �                     @p       q                    �?z�G�z�?             @������������������������       �                      @r       s                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @u       v                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?x                           @�2�tk~�?             "@y       ~       (             �?����>4�?             @z       }                    �?      �?             @{       |                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    �?�XS�_��?Z            �b@�       �                    �?r�q��?;             X@�       �                    �?e�J���?4             U@�       �                    @8����?,            @R@�       �                    @5�_�M"�?            �G@�       �       )             �?����>�?             ?@�       �                    �?n�����?             2@�       �                    @      �?              @������������������������       �                     @������������������������       �                     @�       �                     @���(\��?             $@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?؇���X�?             @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    @�؉�؉�?
             *@�       �                     @���Q��?             @�       �       !             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                     @      �?              @�       �       #             �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    �?      �?	             0@������������������������       �                      @�       �                    �?և���X�?             ,@�       �       !             �?����X�?             @������������������������       �                     @������������������������       �                      @�       �                    �?؇���X�?             @������������������������       �                     �?������������������������       �                     @�       �                     @(ݾ�z��?             :@�       �                    �?�lO���?             3@�       �                    �?�q�q�?             @�       �                    @      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @�       �       
             �?$�q-�?             *@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     "@�       �                    �?����X�?             @������������������������       �                     @������������������������       �                      @�       �                     @������?             &@�       �                     �?      �?             @������������������������       �                      @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?؇���X�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �?�������?             (@�       �                    �?      �?              @������������������������       �                     @������������������������       �                     �?�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?�       �                    @:��\H�?            �J@�       �       %             �?Lh/����?             2@�       �                    @�Q����?             @������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?&�q-�?
             *@�       �       $             �?      �?              @�       �                    @����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                    �?z�G�z�?             @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                    �?VR�s&�?            �A@�       �                    @.�?�P��?             >@�       �                     �?�r����?	             .@�       �                    �?����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                     .@������������������������       �                     @�t�b��     h�h)h,K ��h.��R�(KK�KK��h�B�*       �D@      F@     �S@     @U@     �K@      C@      ;@      ?@     �N@      J@      (@      $@      @      *@      C@      D@      "@      @      �?      "@      ,@      B@      @      @      �?      "@      "@                              �?      "@                                               @                                      �?      �?                                      �?                                                      �?                                                      "@                                              @      B@      @      @                       @      3@              @                       @      3@                                      �?      �?                                      �?                                                      �?                                      �?      2@                                              ,@                                      �?      @                                      �?      �?                                      �?                                                      �?                                              @                                                              @                      @      1@      @                              @      (@      �?                               @      &@                                              @                                       @      @                                              @                                       @                                              �?      �?      �?                                      �?      �?                                              �?                                      �?                                      �?                                                      @      @                                      @      @                                      @      �?                                              �?                                      @                                                      @                                               @              @      @      8@      @       @      �?      @      @                                      @       @                                      @                                                       @                                               @                                                      8@      @       @      �?                      8@      @              �?                      .@                                              "@      @              �?                      @                                              @      @              �?                       @      @              �?                       @                      �?                      �?                      �?                      �?                                                                      �?                      �?                                                      @                                      @                                                               @              5@      2@      7@      (@      @      @      @      @      4@      "@       @      @       @      @      1@      @      �?       @       @      @                                              @                                       @      �?                                      �?      �?                                      �?                                                      �?                                      �?                                                      �?      1@      @      �?       @              �?      0@      �?      �?      �?              �?      0@                                              0@                                      �?                                                              �?      �?      �?                                      �?      �?                                      �?                                                      �?                              �?                                      �?       @              �?                               @                                      �?                      �?                      �?                                                                      �?      �?              @      @      �?       @      �?               @                       @      �?               @                      �?      �?                                      �?      �?                                                                                      �?                       @                                                                      �?                      �?      @      �?                              �?              �?                              �?                                                              �?                                      @                      2@      &@      @      @      �?       @      2@      $@      �?                              0@                                               @      $@      �?                               @       @                                      �?                                              �?       @                                              @                                      �?      @                                               @                                      �?       @                                      �?                                                       @                                               @      �?                                       @                                                      �?                                      �?       @      @      �?       @              �?       @      @      �?                      �?       @              �?                      �?       @                                               @                                      �?                                                                      �?                                      @                                                               @      ,@      *@      2@     �@@     �E@      <@      *@      $@      1@      8@      8@       @      *@      "@      $@      8@      5@      @      $@       @      "@      2@      5@      @      $@       @      "@      1@      @               @       @      "@      .@      @              �?       @      @      @      @                              @              @                              @                                                              @              �?       @      �?      @                               @      �?                                              �?                                       @                                      �?                      @                                              @                      �?                       @                                               @                      �?                                              �?              @      "@                                      @       @                                      �?       @                                      �?                                                       @                                       @                              �?                      @                      �?                      @                                              @                      �?                                                                      @                       @      @               @                                               @                       @      @                                       @      @                                              @                                       @                                              @      �?                                              �?                                      @                                                                      �?      2@      @                              �?      0@       @                                      @       @                                       @       @                                               @                                       @                                               @                                      �?      (@                                      �?      @                                              @                                      �?                                                      "@                                               @      @                                              @                                       @              @      �?      �?      @                      @      �?                                       @                                              �?      �?                                              �?                                      �?                                                              �?      @                                      �?      �?                                              �?                                      �?                                                      @                              �?      @              @      �?                      @                      �?                      @                                                                      �?              �?                      @                                              @                      �?                                      �?      @      �?      "@      3@      4@      �?      @      �?      @      @                      @      �?      �?                              @                                                      �?      �?                                      �?                                                      �?                      �?                      @      @              �?                       @      @                                       @      @                                       @                                                      @              �?                                                                      @      �?                                       @      �?                                       @                                                      �?                                       @                                               @      *@      4@                               @      *@      .@                               @      *@                                       @      @                                              @                                       @                                                       @                                                      .@                                              @�t�bubhhubh)��}�(hhhhhNhKhKhG        hKhNhJC�NhG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKӅ�h��B(.         �       &             �?��2@32�?�            `u@       I       
             �?��ENn�?r            �g@       $                    �?Ӈ0���?9            �X@              !             �?�j;���?            �F@                           �?4և����?	             ,@                           �?      �?             @������������������������       �                      @������������������������       �                      @	                           @{�G�z�?             $@
                           �?r�q��?             @������������������������       �                     @������������������������       �                     �?                           �?      �?             @                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?       !                    �?��_[��?             ?@              	             �?������?             <@                           @      �?             8@                           �?���y4F�?             3@������������������������       �                     $@                           �?X�<ݚ�?             "@������������������������       �                     @              #             �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @              #             �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @               "             �?      �?             @������������������������       �                      @������������������������       �                      @"       #                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @%       4                    @�AMĹ�?             K@&       1                    �?*x9/��?             <@'       0                     @0\�Uo��?
             3@(       /       "             �?0��b�/�?             .@)       .                    �?}��7�?             &@*       -                    �?VUUUUU�?             @+       ,                    @      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @2       3       "             �?�q�q�?             "@������������������������       �                     @������������������������       �                     @5       6                    �?b'vb'v�?             :@������������������������       �                     @7       >                    @�û��|�?             7@8       =                    �?r�q��?             (@9       :       	             �?ףp=
�?             $@������������������������       �                      @;       <                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @?       @                    �?���|���?             &@������������������������       �                     @A       B                    �?      �?              @������������������������       �                     �?C       D                    �?և���X�?             @������������������������       �                     �?E       F                    @      �?             @������������������������       �                      @G       H                      @      �?             @������������������������       �                     �?������������������������       �                     @J       i                    @~<SvL�?9             W@K       d                    �?��>L�*�?            �C@L       [                    �?>��R	�?             ?@M       Z                    �?�q�q�?             8@N       Y                    @�t����?             1@O       X                    �?X�<ݚ�?             "@P       S       #             �?      �?              @Q       R                    @�q�q�?             @������������������������       �                     �?������������������������       �                      @T       W                    �?z�G�z�?             @U       V                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @\       ]                     @����>4�?             @������������������������       �                      @^       c       $             �?�Q����?             @_       `                    �?      �?             @������������������������       �                      @a       b                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?e       h                    �?      �?              @f       g                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @j       y                    �?4uJ0��?            �J@k       p                    @&���^B�?             B@l       m                     �?և���X�?	             ,@������������������������       �                     @n       o       #             �?�q�q�?             "@������������������������       �                     @������������������������       �                     @q       t                    @��!pc�?             6@r       s                     �?���Q��?             @������������������������       �                      @������������������������       �                     @u       v       	             �?�t����?	             1@������������������������       �                     (@w       x       '             �?���Q��?             @������������������������       �                     @������������������������       �                      @z       �                    �?��.k���?	             1@{       �                     �?���!pc�?             &@|       }                    @z�G�z�?             $@������������������������       �                     @~                           �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �?�l�?�d�?f            �b@�       �                    �?,��I�?9            �U@�       �                    �?�r����?             .@������������������������       �        
             *@������������������������       �                      @�       �                    �?�q�q�?.             R@�       �                    �?R=6�z�?(            @P@�       �                    �?��x_F-�?            �I@�       �                    �?��R[s�?            �A@�       �                    �?¦	^_�?             ?@������������������������       �                      @�       �                    �?>���Rp�?             =@�       �                     @r�q��?             8@������������������������       �                     *@�       �                     �?���|���?             &@������������������������       �                     @�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                    �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                    @      �?
             0@������������������������       �                     $@�       �                    �?r�q��?             @������������������������       �                     �?������������������������       �                     @�       �       "             �?X�Cc�?
             ,@�       �                    @�	j*D�?	             *@������������������������       �                      @�       �       )             �?z�G�z�?             @������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                    �?����X�?             @�       �                    �?���Q��?             @������������������������       �                     �?�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    �?     �?-             P@�       �                    @��s��?'            �J@�       �                    �?"���[�?!            �F@�       �       (             �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �       (             �?>��C��?            �E@�       �                    �?¦�F0�?            �D@�       �                    �?      �?              @������������������������       �                      @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     @�       �                    �?�m펠�?            �@@�       �                    �?      �?             @@�       �                    @z�G�z�?             $@������������������������       �                     �?�       �       !             �?�����H�?             "@������������������������       �                     @�       �                    @�q�q�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     6@������������������������       �                     �?������������������������       �                      @�       �                     �?      �?              @������������������������       �                     @�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                     @�C��2(�?             &@������������������������       �                     "@�       �       #             �?      �?              @������������������������       �                     �?������������������������       �                     �?�t�bh�h)h,K ��h.��R�(KK�KK��h�B�'        F@      N@     @R@      S@      O@      ;@      @      @     �A@      M@     �N@      9@      @      @      8@      :@      9@      ,@       @      @      @      3@      @      @       @       @      @      @      �?      �?       @       @                                       @                                                       @                                                      @      @      �?      �?                      @      �?                                      @                                                      �?                                               @      �?      �?                               @      �?                                       @                                                      �?                                                      �?               @      �?      0@      @      @                              0@      @      @                              0@      @      @                              .@              @                              $@                                              @              @                              @                                              �?              @                              �?                                                              @                              �?      @                                      �?                                                      @                                               @       @                                               @                                       @                       @      �?                                              �?                                       @                                       @       @      2@      @      2@      @               @      .@      @       @      @               @      "@      @       @                       @      @      @       @                       @      @       @       @                       @               @       @                       @                       @                       @                                                                       @                                       @                                      @                                                      @                                      @                                              @                      @                      @                                                                      @       @              @      �?      0@      @                      @                               @                      �?      0@      @       @                      �?      "@                                      �?      "@                                               @                                      �?      �?                                      �?                                                      �?               @                                                                              @      @                                      @                                              @      @                                      �?                                              @      @                                              �?                                      @      @                                       @                                              �?      @                                      �?                                                      @       @              &@      @@      B@      &@       @              &@      8@       @               @              @      6@      �?                              @      3@                                      @      (@                                      @      @                                      @      @                                      �?       @                                      �?                                                       @                                      @      �?                                      �?      �?                                              �?                                      �?                                              @                                                      �?                                               @                                              @                       @              �?      @      �?               @                                                              �?      @      �?                                      @      �?                                       @                                              �?      �?                                      �?                                                      �?                              �?                                              @       @      �?                                       @      �?                                       @                                                      �?                              @                                                       @      A@      &@                               @      :@       @                              @       @                                              @                                      @      @                                              @                                      @                                               @      2@       @                               @      @                                       @                                                      @                                              .@       @                                      (@                                              @       @                                      @                                                       @                                       @      "@                                       @      @                                       @       @                                      @                                              @       @                                      @                                                       @                                              �?                                              @      C@      K@      C@      2@      �?       @     �B@      I@                                      *@       @                                      *@                                                       @                                      8@      H@                                      3@      G@                                      $@     �D@                                      "@      :@                                      "@      6@                                       @                                              @      6@                                      @      4@                                              *@                                      @      @                                              @                                      @      �?                                              �?                                      @                                              @       @                                      @                                                       @                                              @                                      �?      .@                                              $@                                      �?      @                                      �?                                                      @                                      "@      @                                      "@      @                                       @                                              �?      @                                              @                                      �?      �?                                              �?                                      �?                                                      �?                                      @       @                                      @       @                                              �?                                      @      �?                                              �?                                      @                                               @                                              �?      @      C@      2@      �?       @      �?      @     �B@       @      �?       @      �?      @      A@      @      �?      �?      �?                                      �?      �?                                                                                      �?              @      A@      @      �?                       @      A@      @      �?                       @      @       @                               @                                                      @       @                                               @                                      @                                              >@       @      �?                              >@       @                                       @       @                                              �?                                       @      �?                                      @                                               @      �?                                      �?      �?                                              �?                                      �?                                              �?                                              6@                                                              �?                       @                                                      @      @              �?                      @                                                      @              �?                                              �?                              @                                      �?      $@                                              "@                                      �?      �?                                              �?                                      �?                        �t�bubhhubh)��}�(hhhhhNhKhKhG        hKhNhJ�R�[hG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKՅ�h��B�.         b       %             �?.��ߴ��?�            `u@                           �?_��}�V�?e            `c@                           �?0�����?
             ,@                           �?r�q��?	             (@������������������������       �                     $@������������������������       �                      @������������������������       �                      @       O                    �?}�)��?[            �a@	       0                    @�Jup��?D            �Z@
       +                    @�Cc}h��?%             L@       $                    �?o�`� �?!            �I@                           �?$��,�?            �E@                           �?$I�$I��?
             ,@                           @0�����?             @              (             �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?                           �?�$I�$I�?             @                           @�q�q�?             @                           �?z�G�z�?             @������������������������       �                      @              (             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     �?       #                    �?�-Z�?             =@       "                    �?@4և���?             <@       !                    �?�t����?
             1@               "             �?      �?              @������������������������       �                     @������������������������       �                      @������������������������       �                     "@������������������������       �                     &@������������������������       �                     �?%       &       '             �?      �?              @������������������������       �                     @'       *                    �?      �?             @(       )                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @,       /       	             �?z�G�z�?             @-       .                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @1       @                    �?|�/L�
�?             I@2       ?                    �?����>�?             <@3       8                    @���B���?             :@4       7                    �?H�z�G�?             $@5       6                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @9       <                     �?      �?
             0@:       ;                    @$�q-�?             *@������������������������       �                     (@������������������������       �                     �?=       >                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @A       N                    �?n,�Ra�?             6@B       G                    �?�G�z��?             4@C       D                    �?      �?              @������������������������       �                     @E       F       #             �?      �?              @������������������������       �                     �?������������������������       �                     �?H       M       !             �?r�q��?             (@I       J                     @�C��2(�?             &@������������������������       �                      @K       L                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @P       _                    �?PuPu�?            �A@Q       R       )             �?7�ٔ_�?             =@������������������������       �                     .@S       T                    �?������?             ,@������������������������       �                      @U       ^       $             �?�q�q�?	             (@V       Y                    �?2(&ޏ�?             &@W       X                    @      �?              @������������������������       �                     �?������������������������       �                     �?Z       [                    �?�����H�?             "@������������������������       �                     @\       ]                     @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?`       a                    @      �?             @������������������������       �                     @������������������������       �                     @c       �                    �?��a��*�?r            `g@d       �                    @)+#��?h            `e@e       �                    @$�/�߹�?Q            �a@f       �                    @���Q��?8            @X@g       z                    @�����Y�?/             T@h       u                    �?� u#��?             C@i       r       $             �?      �?             @@j       m                    �?      �?
             4@k       l                    �?�8��8��?             (@������������������������       �                     �?������������������������       �                     &@n       o                    �?      �?              @������������������������       �                     @p       q                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @s       t                    @�8��8��?             (@������������������������       �                     &@������������������������       �                     �?v       w                    �?�q�q�?             @������������������������       �                     @x       y                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @{       �                    �?������?             E@|       �                    �?     ��?             @@}       �                    �?��S�r
�?             <@~       �                    �?��ջ���?             :@       �                    �?��8��8�?	             (@�       �                    �?      �?              @������������������������       �                      @������������������������       �                     @�       �                    �?      �?             @������������������������       �                      @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?�m۶m��?	             ,@������������������������       �                     "@�       �                    �?{�G�z�?             @�       �                    �?�q�q�?             @������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    @p=
ףp�?             $@�       �                    �?      �?              @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    @�M�]��?	             1@�       �                    �?����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     $@�       �       
             �?��ճC��?             F@�       �                    @(������?             3@������������������������       �                     ,@�       �       !             �?���Q��?             @������������������������       �                     @������������������������       �                      @�       �                    �?�l�����?             9@�       �                    �?�mM`���?             7@�       �                    �?|�/��>�?             1@�       �       '             �?�8��8��?             (@�       �                    @r�q��?             @������������������������       �                     @�       �       #             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �?{�G�z�?             @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                      @�       �                    �?���ĳ��?             >@�       �                    @���!pc�?             &@������������������������       �                      @������������������������       �                     @�       �                    �?��|���?             3@�       �                    @f�t���?             1@�       �                    �?�<ݚ�?             "@������������������������       �                     �?�       �                    �?      �?              @�       �       #             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �       !             �?      �?              @������������������������       �                     @�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    �?     ��?
             0@�       �                    �?�	j*D�?             *@�       �                     @"pc�
�?             &@�       �                    �?      �?              @������������������������       �                     @������������������������       �                     �?�       �       #             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @�t�bh�h)h,K ��h.��R�(KK�KK��h�B�'        >@     �L@     @V@     @U@     �L@      8@      =@      L@      G@      4@      �?      @      $@       @                               @      $@                                       @      $@                                                                                       @               @                                      3@      K@      G@      4@      �?      �?      2@     �G@      7@      0@      �?      �?      1@     �@@      @              �?              *@      @@      @              �?               @      ?@      @              �?              @      @      @                              @      �?      �?                              @      �?                                      @                                                      �?                                                      �?                              �?      @       @                                      @       @                                      @      �?                                       @                                               @      �?                                              �?                                       @                                                      �?                              �?                                               @      :@                      �?               @      :@                                       @      .@                                       @      @                                              @                                       @                                                      "@                                              &@                                                                      �?              @      �?       @                              @                                              �?      �?       @                              �?      �?                                      �?                                                      �?                                                       @                              @      �?                                      �?      �?                                              �?                                      �?                                              @                                              �?      ,@      2@      0@              �?      �?      @      "@      ,@              �?      �?      @      @      ,@              �?      �?      @      @                              �?      @                                              @                                      �?                                                              @                                              �?      ,@              �?                              (@              �?                              (@                                                              �?                      �?       @                                      �?                                                       @                                       @                                      &@      "@       @                              &@      "@                                      �?      @                                              @                                      �?      �?                                              �?                                      �?                                              $@       @                                      $@      �?                                       @                                               @      �?                                       @                                                      �?                                              �?                                                       @                      �?      @      7@      @                      �?      @      7@      �?                                      .@                              �?      @       @      �?                               @                                      �?       @       @      �?                      �?      �?       @      �?                      �?      �?                                      �?                                                      �?                                                       @      �?                                      @                                              @      �?                                      @                                                      �?                              �?                                              @              @                              @                                                              @                      �?      �?     �E@     @P@      L@      5@      �?      �?      A@      O@      L@      1@      �?      �?      A@      N@      D@      @              �?      @@     �B@      8@      @              �?      >@      @@      ,@      @              �?      <@      "@                              �?      :@      @                                      .@      @                                      &@      �?                                              �?                                      &@                                              @      @                                      @                                              �?      @                                      �?                                                      @                              �?      &@                                              &@                                      �?                                                       @      @                                              @                                       @      �?                                              �?                                       @                                               @      7@      ,@      @                       @      0@      *@      �?                       @      0@      "@      �?                      �?      0@       @      �?                              @      @      �?                               @      @                                       @                                                      @                                      @              �?                               @                                              �?              �?                              �?                                                              �?                      �?      &@       @                                      "@                                      �?       @       @                              �?               @                                              �?                              �?              �?                              �?                                                              �?                                       @                                      �?              �?                              �?                                                              �?                                              @                                      @      �?       @                              @      �?                                      �?      �?                                      �?                                                      �?                                      @                                                               @                       @      @      $@                               @      @                                              @                                       @                                                              $@              �?               @      7@      0@       @                              ,@      @       @                              ,@                                                      @       @                                      @                                                       @      �?               @      "@      *@              �?               @      @      *@              �?               @      �?      *@                                      �?      &@                                      �?      @                                              @                                      �?       @                                               @                                      �?                                                      @              �?               @               @              �?                               @              �?                                                                               @                               @                                                      @                                               @                                               @      0@      (@                                       @      @                                       @                                                      @                               @       @      "@                               @       @      @                               @      @                                      �?                                              �?      @                                      �?       @                                      �?                                                       @                                              @                                              �?      @                                              @                                      �?      @                                      �?                                                      @                                               @                      "@      @              @                      "@                      @                      "@                       @                      @                      �?                      @                                                                      �?                       @                      �?                                              �?                       @                                                                       @                              @                �t�bubhhubh)��}�(hhhhhNhKhKhG        hKhNhJ�v}hG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK���h��B8*         �                    @���ܨ��?�            `u@       [                    �?�_�3lF�?�            @s@                           �?�c�,:#�?_            �b@                           �?���>*�?            �C@������������������������       �                     .@                           �?��8��8�?             8@              #             �?�q�q�?             (@                            @�$I�$I�?             @	       
       &             �?z�G�z�?             @������������������������       �                     @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                           �?���Q��?             @                           @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @                           �?�8��8��?             (@                           @      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     @       $                    �?PE=l18�?H            �[@       !                    �?      �?             (@              '             �?      �?              @������������������������       �                      @                             @      �?             @              %             �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?"       #                      @      �?             @������������������������       �                     @������������������������       �                     �?%       B       &             �?�����?@            �X@&       ;                    �?���Y �?             ;@'       :                    @ףp=
��?             4@(       9                    �?��ӭ�a�?             2@)       0                    �?���Er�?             1@*       /                    �?{�G�z�?             @+       ,                    �?�q�q�?             @������������������������       �                     �?-       .                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @1       8                    �?      �?             (@2       3                    �?"pc�
�?             &@������������������������       �                     @4       7                    @      �?              @5       6                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @<       ?                    �?�$I�$I�?             @=       >                    @z�G�z�?             @������������������������       �                     @������������������������       �                     �?@       A                    �?      �?              @������������������������       �                     �?������������������������       �                     �?C       R                    �?"赢<6�?-            �Q@D       M                    �?"pc�
�?             F@E       F                    �?������?            �B@������������������������       �                     9@G       H                    �?�q�q�?             (@������������������������       �                     @I       L                    �?      �?              @J       K       $             �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @N       O       '             �?և���X�?             @������������������������       �                     @P       Q       !             �?      �?             @������������������������       �                     �?������������������������       �                     @S       X       
             �?���^�?             ;@T       U                    �?���}<S�?             7@������������������������       �                     2@V       W       !             �?���Q��?             @������������������������       �                     @������������������������       �                      @Y       Z                    �?      �?             @������������������������       �                     �?������������������������       �                     @\       �                    @<�1�'��?\            �c@]       �       %             �?�l'l��?F             _@^                           �?u{H���?'            @Q@_       j       #             �?J]�'GZ�?            �G@`       g       
             �?�^B{	��?             2@a       f                    �?:/����?             ,@b       e       	             �?�g���e�?             &@c       d                    �?�z�G��?             $@������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     @h       i                    �?      �?             @������������������������       �                     �?������������������������       �                     @k       |                    �?��л��?             =@l       {                    �?2U0*��?             9@m       r                    �?r�q��?             8@n       o                    �?      �?             @������������������������       �                      @p       q                    �?      �?              @������������������������       �                     �?������������������������       �                     �?s       t                    @R���Q�?
             4@������������������������       �                     $@u       x                     @�z�G��?             $@v       w                    @z�G�z�?             @������������������������       �                     @������������������������       �                     �?y       z                    �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?}       ~                    @      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �?�i�V��?
             6@�       �       $             �?�\��N��?	             3@�       �       !             �?؇���X�?             ,@������������������������       �                     (@������������������������       �                      @�       �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    �?
ףp=
�?            �K@�       �                    @ޯ�f��?             C@�       �                    �?~h����?             <@�       �                    �?H�z�G�?             4@������������������������       �                      @�       �                    �?�q�q�?             2@�       �       "             �?8�Z$���?	             *@�       �                    �?�8��8��?             (@������������������������       �                      @�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �                    �?z�G�z�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    �?ףp=
�?             $@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    �?�M�]��?             1@������������������������       �                      @�       �                    �?�����H�?             "@������������������������       �                     �?������������������������       �                      @�       �                    �?4��g�?            �A@�       �                    @�t��q3�?             =@�       �                    �?8��8���?             8@�       �                    @�KM�]�?
             3@�       �                    �?z�G�z�?             $@������������������������       �                     @�       �                    @���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     "@�       �                    �?�Q����?             @�       �                    �?      �?             @������������������������       �                      @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    @��\���?             A@�       �                    �?�KM�]�?             3@�       �                    @�X�<ݺ?             2@������������������������       �                     �?������������������������       �                     1@������������������������       �                     �?�       �                    �?z�G�z�?	             .@������������������������       �                     (@������������������������       �                     @�t�b��#     h�h)h,K ��h.��R�(KK�KK��h�B0$        B@     @P@     @T@     @U@      G@      =@      B@     @P@     @T@     �T@      :@      1@      :@      D@      F@      2@      (@      "@      1@      �?      ,@               @      @      .@                                               @      �?      ,@               @      @       @      �?      @               @      @       @      �?                              @              �?                              @                                              @              �?                              �?              �?                                                                              �?       @                                                              @               @                              �?               @                              �?                                                               @                               @                                              &@                      �?                      @                      �?                      @                                                                      �?                      @                              "@     �C@      >@      2@      $@      @      �?              �?      @      @      @      �?              �?      @               @                                               @      �?              �?      @                                      �?      @                                      �?                                                      @                      �?                                                                              @      �?                                      @                                                      �?       @     �C@      =@      ,@      @      �?              @      @      &@      @      �?               @      @      &@      �?      �?                      @      &@      �?      �?                      @      &@      �?                               @       @      �?                               @              �?                              �?                                              �?              �?                                              �?                              �?                                                       @                                      @      "@                                       @      "@                                              @                                       @      @                                       @       @                                               @                                       @                                                      @                                      �?                                                                      �?               @                                              �?       @              @                              �?              @                                              @                              �?                                      �?      �?                                      �?                                                      �?                               @      B@      6@      @       @               @      B@                                      @     �@@                                              9@                                      @       @                                              @                                      @      @                                      @      �?                                      @                                                      �?                                              @                                      @      @                                      @                                              �?      @                                      �?                                                      @                                                      6@      @       @                              5@               @                              2@                                              @               @                              @                                                               @                              �?      @                                      �?                                                      @                      $@      9@     �B@     @P@      ,@       @      "@      7@      B@     �C@      "@       @      @      7@      7@      0@                      @      &@      7@      @                      �?      @      @      @                      �?      @      @      @                      �?      @      @                                      @      @                                              @                                      @                                      �?                                                                      @                                      @      �?                                              �?                                      @                              @      @      1@      @                       @      @      1@      @                      �?      @      1@      @                      �?      @                                               @                                      �?      �?                                      �?                                                      �?                                                      1@      @                                      $@                                              @      @                                      @      �?                                      @                                                      �?                                      @       @                                      @                                                       @                      �?                                              @      �?                                      @                                                      �?                                      �?      (@              "@                      �?      (@              @                              (@               @                              (@                                                               @                      �?                      @                                              @                      �?                                                                      @                       @              *@      7@      "@       @       @              (@      .@      "@               @              (@      ,@                       @              (@      @                       @                                                              (@      @                                      &@       @                                      &@      �?                                       @                                              @      �?                                      @                                                      �?                                              �?                                      �?      @                                      �?      �?                                      �?                                                      �?                                              @                                               @                                              �?      "@                                      �?      �?                                      �?                                                      �?                                               @                              �?       @               @                               @                                      �?                       @                      �?                                                                       @      �?       @      �?      :@      @              �?       @      �?      4@      @              �?       @      �?      4@                               @              1@                               @               @                                              @                               @              @                               @                                                              @                                              "@                      �?              �?      @                      �?                      @                                               @                      �?                      �?                                              �?                      �?                                                              �?                                                              @                                      @                                               @      4@      (@                               @      1@                                      �?      1@                                      �?                                                      1@                                      �?                                                      @      (@                                              (@                                      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hKhNhJg}�XhG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK���h��Bx(         0                    �?�p���?�            `u@       !                     �?�o+��?>            �W@       
                    �?      �?*             P@                           @�	j*D�?	             *@������������������������       �                     @                           �?և���X�?             @������������������������       �                     @       	                    �?      �?             @������������������������       �                     @������������������������       �                     �?               !             �?�t����?!            �I@                           @      �?             D@                           �?�S����?             3@������������������������       �                     "@                           �?�z�G��?             $@������������������������       �                     @                           �?      �?             @������������������������       �                     �?              #             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?                           �?և���X�?             5@                           @���Q��?             .@                           �?      �?             (@������������������������       �                     @              $             �?      �?             @                           �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �        
             &@"       '                    �?�P�*�?             ?@#       &       '             �?      �?	             0@$       %       $             �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     (@(       -                    �?z�G�z�?             .@)       ,                    �?�8��8��?	             (@*       +                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@.       /       #             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?1       �       &             �?ho*ϕj�?�            �n@2       [                    @ \�F�)�?i            �c@3       T       "             �?���l<�?4            @S@4       G                    @     t�?+             P@5       B                    �?�99lMt�?            �C@6       ?                    �?�-Z�?             =@7       8                    @�6|����?             :@������������������������       �        	             1@9       >                    �?h/�����?             "@:       ;                    �?�$I�$I�?             @������������������������       �                      @<       =                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @@       A       !             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @C       F       )             �?���Q��?             $@D       E                     �?      �?              @������������������������       �                      @������������������������       �                     @������������������������       �                      @H       M                    �? �o_��?             9@I       L                    �?      �?
             0@J       K                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     $@N       O                    �?�q�q�?             "@������������������������       �                     @P       Q                    �?      �?             @������������������������       �                      @R       S       )             �?      �?              @������������������������       �                     �?������������������������       �                     �?U       Z                      @$�q-�?	             *@V       Y                    �?      �?             @W       X                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     "@\       �                    �?H�z��?5             T@]       r                    @�OY>{�?-            @P@^       i                    �?�8��8��?             8@_       h                    �?��S���?
             .@`       g                    �?/����?	             ,@a       f       $             �?������?             @b       c       )             �?      �?             @������������������������       �                      @d       e                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?j       k       #             �?h/�����?             "@������������������������       �                      @l       q                    �?�$I�$I�?             @m       p                    �?�q�q�?             @n       o                    �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?s       �                     @��r._�?            �D@t       u                    �?�C��2(�?            �@@������������������������       �        	             *@v       {                    �?R���Q�?             4@w       z                    �?@4և���?	             ,@x       y                    �?r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @|       }                    �?�q�q�?             @������������������������       �                     �?~                           �?z�G�z�?             @������������������������       �                     �?�       �                     @      �?             @������������������������       �                     @������������������������       �                     �?�       �                    @      �?              @������������������������       �                     @������������������������       �                     @�       �                    �?z�G�z�?             .@������������������������       �                     &@�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �?��a���?4            �V@�       �                    �?6�h$��?            �F@������������������������       �        
             2@�       �                    �?��E���?             ;@�       �                    �?
ףp=
�?             $@�       �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    �?�Q����?             @������������������������       �                     �?�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �?�t����?             1@�       �       '             �?�eP*L��?             &@������������������������       �                      @�       �                    �?�q�q�?             "@�       �                    @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �       #             �??7(�Q�?            �F@�       �                    �?������?             1@�       �                    �?      �?              @�       �       $             �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     "@�       �                    @      �?             <@�       �                    �?h/�����?             2@�       �       )             �?�z�G��?             $@������������������������       �                     @�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �?      �?              @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?z�G�z�?             @�       �                    @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     $@�t�bh�h)h,K ��h.��R�(KK�KK��h�B�"        G@     �N@      V@      R@      K@      5@      E@     �J@                                      8@      D@                                      "@      @                                      @                                              @      @                                              @                                      @      �?                                      @                                                      �?                                      .@      B@                                      .@      9@                                      @      0@                                              "@                                      @      @                                              @                                      @      �?                                      �?                                               @      �?                                       @                                                      �?                                      (@      "@                                      @      "@                                      @      "@                                              @                                      @      @                                      �?      @                                      �?                                                      @                                       @                                              @                                              @                                                      &@                                      2@      *@                                      .@      �?                                      @      �?                                              �?                                      @                                              (@                                              @      (@                                      �?      &@                                      �?      �?                                      �?                                                      �?                                              $@                                       @      �?                                       @                                                      �?                                      @       @      V@      R@      K@      5@                      A@     �H@     �J@      5@                      A@      E@      �?                             �@@      >@      �?                              :@      (@      �?                              6@      @      �?                              5@      @      �?                              1@                                              @      @      �?                               @      @      �?                               @                                                      @      �?                                      @                                                      �?                               @                                              �?       @                                      �?                                                       @                                      @      @                                       @      @                                       @                                                      @                                       @                                              @      2@                                      �?      .@                                      �?      @                                              @                                      �?                                                      $@                                      @      @                                      @                                              �?      @                                               @                                      �?      �?                                              �?                                      �?                                              �?      (@                                      �?      @                                      �?      �?                                              �?                                      �?                                                       @                                              "@                                              @      J@      5@                              @      D@      2@                              @      @      &@                              @       @      $@                              @      �?      $@                              @      �?      @                              @      �?                                       @                                              �?      �?                                              �?                                      �?                                                              @                                              @                                      �?                                      @      @      �?                               @                                               @      @      �?                               @      @                                       @      @                                       @                                                      @                                              �?                                                      �?                                      A@      @                                      >@      @                                      *@                                              1@      @                                      *@      �?                                      @      �?                                              �?                                      @                                               @                                              @       @                                              �?                                      @      �?                                      �?                                              @      �?                                      @                                                      �?                                      @      @                                      @                                                      @                                      (@      @                                      &@                                              �?      @                                      �?                                                      @      @       @      K@      7@      �?              @      @     �@@      �?      �?                              2@                              @      @      .@      �?      �?              @      �?      @      �?      �?              @      �?                                      @                                                      �?                                                      @      �?      �?                                              �?                              @      �?                                      @                                                      �?                              @      (@                                      @      @                                       @                                              @      @                                      @      �?                                      @                                                      �?                                              @                                              @                                       @      5@      6@                                      *@      @                                      @      @                                      @      �?                                              �?                                      @                                                      @                                      "@                                       @       @      2@                               @       @       @                                      @      @                                      @                                              �?      @                                              @                                      �?                                       @      �?      @                               @              �?                                              �?                               @                                                      �?      @                                      �?       @                                      �?                                                       @                                               @                                              $@                �t�bubhhubh)��}�(hhhhhNhKhKhG        hKhNhJ	�tlhG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKۅ�h��B�/         |       
             �?n	#N;��?�            `u@       A       %             �?C�Im_�?{            �h@       "                     @��~����?E            @\@                           �?�U����?            �H@������������������������       �                     @              "             �?��J��?             F@                           @>��R	�?             ?@              !             �?H��	,U�?             7@	                           �?��!pc�?             &@
                           �?      �?              @                           �?�q�q�?             @������������������������       �                     �?                           �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @                           �?�8��8��?             (@������������������������       �                      @                           �?      �?             @������������������������       �                     @������������������������       �                     �?                           �?      �?              @������������������������       �                     �?                           @؇���X�?             @������������������������       �                     @������������������������       �                     �?       !                    �?8�Z$���?             *@                            @�8��8��?             (@                           @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     "@������������������������       �                     �?#       2                    �?     p�?'             P@$       )                    �?��
P��?            �A@%       &       !             �?�����H�?             2@������������������������       �                     $@'       (       "             �?      �?              @������������������������       �                      @������������������������       �                     @*       /                    �?�t����?             1@+       ,       '             �?��S�ۿ?             .@������������������������       �                     "@-       .                    �?r�q��?             @������������������������       �                     �?������������������������       �                     @0       1                    �?      �?              @������������������������       �                     �?������������������������       �                     �?3       @                    @�S�����?             =@4       =                    �?�K8��?             :@5       <       (             �?�8��8��?             8@6       7                     �?�nkK�?             7@������������������������       �                     .@8       ;                    �?      �?              @9       :                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?>       ?                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @B       s                    �?q�9��?6            �T@C       p                    �?^@l*9�?/            �Q@D       ]                    �?*��|6��?)             M@E       V                    �?����>�?             <@F       U                    �?�z�G��?             4@G       P                    @n�����?             2@H       M       $             �?��1G���?	             *@I       L                     �?X�<ݚ�?             "@J       K                    �?؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @N       O                    �?      �?             @������������������������       �                      @������������������������       �                      @Q       T                    �?z�G�z�?             @R       S                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @W       \                    �?      �?              @X       [                    �?      �?             @Y       Z                     �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @^       k                    @�A��S�?             >@_       j                    @d}h���?	             ,@`       a       #             �?t�E]t�?             &@������������������������       �                      @b       i                    �?B{	�%��?             "@c       h                    �?      �?              @d       e                    �?�q�q�?             @������������������������       �                     �?f       g                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @l       o                    @     ��?             0@m       n                    �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �        
             &@q       r       )             �?      �?             (@������������������������       �                     "@������������������������       �                     @t       u                    @g\�5�?             *@������������������������       �                     @v       {                    �?      �?              @w       x                    �?      �?             @������������������������       �                      @y       z                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @}       �                    �?��␸��?[            @b@~       �                    �?�6c���?V             a@       �       %             �?8���:�?G            �[@�       �                    �?(����?            �E@�       �                    �?D�n�3�?             3@�       �                    �?�q�q�?             "@������������������������       �                     @������������������������       �                     @�       �                    �?z�G�z�?             $@�       �       #             �?�����H�?             "@������������������������       �                     @�       �                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                    �?      �?             8@�       �                     @      �?             4@������������������������       �                     @�       �                    �?X�Cc�?             ,@�       �                    @"pc�
�?             &@�       �                    @�q�q�?             @������������������������       �                     @�       �       )             �?�q�q�?             @�       �                     @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �       $             �?�9߄*�?)             Q@�       �                    �?�0��?!             K@�       �                    @��|���?             C@�       �                    @f�t���?             A@�       �                    �?���y4F�?             3@�       �                     @؇���X�?
             ,@������������������������       �                     $@�       �                     �?      �?             @�       �                    �?�q�q�?             @�       �       #             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �       '             �?���Q��?             @������������������������       �                     @������������������������       �                      @�       �                    �?��S�ۿ?             .@������������������������       �        	             *@�       �       #             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    @     ��?	             0@�       �                    @ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     @�       �                    �?/����?             ,@�       �                    @޾�z�<�?             *@������������������������       �                      @�       �       '             �?�C��2(�?             &@������������������������       �                      @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                     @���Mb�?             9@�       �                    �?����X�?             @������������������������       �                     @������������������������       �                      @�       �                    �?�8��8��?             2@�       �                    �?0�����?             ,@�       �                     @�$I�$I�?             @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �?؇���X�?             @������������������������       �                     @������������������������       �                     �?�       �                    @      �?             @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                    �?p=
ףp�?             $@�       �                     �?�<ݚ�?             "@������������������������       �                     @�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?�t�bh�h)h,K ��h.��R�(KK�KK��h�B)       �J@     �P@     �R@      T@      L@      (@     �C@     �I@      I@      ?@      2@      @      A@      G@      <@       @              @      0@      ;@      @      �?                      @                                              &@      ;@      @      �?                      &@      0@      @      �?                      @      .@      @                              @      @       @                               @      @       @                                      @       @                                              �?                                      @      �?                                              �?                                      @                                       @                                              @                                                      &@      �?                                       @                                              @      �?                                      @                                                      �?                              @      �?              �?                                              �?                      @      �?                                      @                                                      �?                                              &@       @                                      &@      �?                                       @      �?                                              �?                                       @                                              "@                                                      �?                              2@      3@      7@      �?              @      2@      1@                                      0@       @                                      $@                                              @       @                                               @                                      @                                               @      .@                                      �?      ,@                                              "@                                      �?      @                                      �?                                                      @                                      �?      �?                                              �?                                      �?                                                       @      7@      �?              @               @      7@      �?                               @      6@                                      �?      6@                                              .@                                      �?      @                                      �?       @                                               @                                      �?                                                      @                                      �?                                                      �?      �?                                              �?                                      �?                                                                      @      @      @      6@      =@      2@      @      @      �?      0@      ;@      2@      @      @      �?      *@      2@      2@      @       @              @      .@      @      �?       @              @       @      @      �?       @              @      @      @      �?       @              @      @       @                              �?      @       @                              �?      @                                      �?                                                      @                                                       @               @               @                                               @                               @                                                                              @      �?                                      @      �?                                      @                                                      �?                                      �?                                       @                                              @      �?                                      @      �?                                      �?      �?                                              �?                                      �?                                               @                                              @                      @      �?      $@      @      &@       @      @      �?      @      �?               @              �?      @      �?               @                                               @              �?      @      �?                                      @      �?                                       @      �?                                      �?                                              �?      �?                                      �?                                                      �?                                      @                                      �?                                      @                                                              @       @      &@                              @       @                                      @                                                       @                                                      &@                              @      "@                                              "@                                      @                                      @      @       @              �?                      @                                      @      �?       @              �?                      �?       @              �?                               @                                      �?                      �?                      �?                                                                      �?              @                                      ,@      .@      9@     �H@      C@      @      *@      *@      9@      E@      C@      @      &@       @      8@      C@      <@       @      &@       @      .@      "@                      &@       @                                      @      @                                              @                                      @                                               @       @                                       @      �?                                      @                                               @      �?                                       @                                                      �?                                              �?                                                      .@      "@                                      .@      @                                      @                                              "@      @                                      "@       @                                      @       @                                      @                                              �?       @                                      �?      �?                                      �?                                                      �?                                              �?                                      @                                                      @                                              @                                      "@      =@      <@       @                      @      =@      2@      �?                      @      0@      2@                              @      0@      ,@                              @      .@                                       @      (@                                              $@                                       @       @                                       @      �?                                      �?      �?                                              �?                                      �?                                              �?                                                      �?                                       @      @                                              @                                       @                                                      �?      ,@                                              *@                                      �?      �?                                              �?                                      �?                                                      @                               @      *@              �?                              "@              �?                              "@                                                              �?                       @      @                                       @                                                      @                                      @              $@      �?                       @              $@      �?                       @                                                              $@      �?                                       @                                               @      �?                                              �?                                       @                              �?                               @      @      �?      @      $@      @       @      @                                              @                                       @                                                              �?      @      $@      @                               @      $@       @                              �?      @       @                              �?               @                                               @                              �?                                                      @                                      �?      @                                              @                                      �?                                      �?       @              �?                      �?       @                                               @                                      �?                                                                      �?      �?       @              @                               @              @                                              @                               @               @                                               @                               @                                      �?                                        �t�bubhhubh)��}�(hhhhhNhKhKhG        hKhNhJ�ޡhG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKׅ�h��B/         �                    �?������?�            `u@                           �?B��︤�?�            �l@                           �?�ɜoB�?             A@              &             �?��Wϊ�?             >@                           @�θ�?	             *@                           @h/�����?             "@       
                    �?z�G�z�?             @       	                      @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     @                           �?�W��H��?             1@                           �?��S�ۿ?	             .@������������������������       �                     ,@������������������������       �                     �?                           �?      �?              @������������������������       �                     �?������������������������       �                     �?                           @      �?             @������������������������       �                     @������������������������       �                     �?       i                    @;j5r��?x            `h@       X                    @��D���?R            @`@       7                    �?ٰ�K2��?<            �W@       (       &             �?�s���?$            �M@                           �?��{ ��?             7@                           @      �?              @������������������������       �                     �?������������������������       �                     @        !                    �?���Q��?             .@������������������������       �                     @"       #                    @      �?              @������������������������       �                     �?$       %                    �?؇���X�?             @������������������������       �                      @&       '       !             �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @)       .                    �?x�5?,R�?             B@*       +                    �?��S�ۿ?             .@������������������������       �        	             (@,       -       	             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?/       0       '             �?AA�?             5@������������������������       �                      @1       6       
             �?޾�z�<�?             *@2       5                     @      �?             @3       4                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     "@8       ?                    �?�n~��?            �A@9       >                    �?�$I�$I�?             @:       ;                     �?�q�q�?             @������������������������       �                     @<       =                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?@       U       !             �?x9/���?             <@A       T                    �?袋.���?             6@B       Q                    �?mdk����?             5@C       P                    �?�q�q�?             2@D       O                    �?      �?	             0@E       L                    �?����X�?             ,@F       K       &             �?�����H�?             "@G       J                    �?؇���X�?             @H       I                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @M       N       '             �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                      @R       S                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?V       W                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?Y       Z                    �?ԭ�a�2�?             B@������������������������       �        	             0@[       f                    �?���Q��?             4@\       a       	             �?�[��"e�?             2@]       `                    @ףp=
�?             $@^       _                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @b       e                    �?      �?              @c       d       '             �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @g       h       '             �?      �?              @������������������������       �                     �?������������������������       �                     �?j       }                    @���#�%�?&            @P@k       p       #             �?:ɨ��?            �@@l       m                    �?      �?	             0@������������������������       �                     *@n       o                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?q       x                    �?@�0�!��?
             1@r       w                    �?���Q��?             $@s       v                    �?և���X�?             @t       u                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @y       |                    �?����X�?             @z       {                     @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @~                           @      �?             @@������������������������       �                      @�       �                    �?�q�q�?             >@�       �       %             �?�n_Y�K�?             :@������������������������       �                     �?�       �                    �?���Q��?             9@�       �       
             �?�eP*L��?	             &@�       �                    @r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    @z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                    @����X�?             ,@������������������������       �                     @������������������������       �                     $@������������������������       �                     @�       �                    �?��j8B9�?H            @\@�       �                    �?��+��?            �B@�       �                     @��Q��?             4@������������������������       �                     (@�       �                     �?      �?              @�       �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    �?ҳ�wY;�?
             1@������������������������       �                     @�       �                    �?���Q��?             $@�       �                     �?؇���X�?             @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                     �?Xp���?2             S@�       �                    @VUUUUU�?             5@�       �                    @8�Z$���?
             *@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?�       �       #             �?�����H�?             "@�       �       '             �?z�G�z�?             @������������������������       �                     @�       �                     �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �       %             �?      �?              @������������������������       �                     �?������������������������       �                     @�       �                    @�*�R�Z�?$            �K@�       �                    �?��)f���?!            �I@�       �                    �?(\���(�?             D@�       �                    @�m펠�?            �@@�       �                     @"pc�
�?             &@������������������������       �                     "@������������������������       �                      @�       �                    �?���7�?             6@�       �                    �?��S�ۿ?	             .@������������������������       �                     &@�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �       !             �?������?             @�       �       (             �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?{�G�z�?             @�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?�       �                    �?"pc�
�?             &@�       �       $             �?X�<ݚ�?             "@�       �                     @z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    �?      �?             @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                    �?      �?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�t�bh�h)h,K ��h.��R�(KK�KK��h�BP(       �C@     �H@      V@     �U@      I@      =@      5@      8@      G@     �Q@      D@      <@      ,@       @      @      @      @      @      ,@       @      @              @      @              �?      @              @      @              �?      @              @                      �?      @                                      �?       @                                      �?                                                       @                                               @                                                              @                                                      @      ,@      �?      �?                      �?      ,@      �?                                      ,@                                                      �?                                                      �?                      �?                      �?                                                                      �?                              @              �?                              @                                                              �?      @      6@     �D@     �P@      B@      6@      @      6@     �D@      N@                      @      4@      C@      @@                      �?      0@      ;@      .@                              �?      "@      *@                              �?              @                              �?                                                              @                                      "@      @                                      @                                               @      @                                      �?                                              �?      @                                               @                                      �?      @                                      �?                                                      @                      �?      .@      2@       @                      �?      ,@                                              (@                                      �?       @                                               @                                      �?                                                      �?      2@       @                                       @                                      �?      $@       @                              �?      �?       @                              �?      �?                                              �?                                      �?                                                               @                                      "@                              @      @      &@      1@                      �?       @      @                                       @      @                                              @                                       @      �?                                       @                                                      �?                              �?                                               @       @      @      1@                      �?       @      @      (@                               @      @      (@                                      @      (@                                      @      $@                                      @      $@                                      �?       @                                      �?      @                                      �?      @                                      �?                                                      @                                              @                                               @                                      @       @                                      @                                                       @                                       @                                                       @                               @      �?                                              �?                                       @                                      �?                                              �?                      @                                              @                      �?                                              @       @      @      <@                                              0@                      @       @      @      (@                      @      �?       @      (@                              �?              "@                              �?              @                                              @                              �?                                                              @                      @               @      @                                       @      @                                       @                                                      @                      @                                                      �?      �?                                              �?                                      �?                                                              @      B@      6@                              @      8@       @                              �?      .@                                              *@                                      �?       @                                               @                                      �?                                              @      "@       @                              @      @                                      @      @                                      @      �?                                      @                                                      �?                                              @                                      @                                                      @       @                                      �?       @                                               @                                      �?                                              @                                              (@      4@                                       @                                              $@      4@                                      $@      0@                                              �?                                      $@      .@                                      @      @                                      @      �?                                      @                                                      �?                                      �?      @                                      �?                                                      @                                      @      $@                                      @                                                      $@                                              @      2@      9@      E@      1@      $@      �?      2@      3@                                      @      *@                                              (@                                      @      �?                                      @      �?                                      @                                                      �?                                      @                                              &@      @                                      @                                              @      @                                      �?      @                                      �?       @                                      �?                                                       @                                              @                                      @                                                      @      E@      1@      $@      �?              �?      @      "@      @                      �?      @       @                              �?      @                                              @                                      �?                                                      �?       @                                      �?      @                                              @                                      �?      �?                                      �?                                                      �?                                              @                                              �?      @                                      �?                                                      @                      @      C@       @      @      �?              @      C@      @       @                      @      @@      @       @                       @      >@      �?                               @      "@                                              "@                                       @                                                      5@      �?                                      ,@      �?                                      &@                                              @      �?                                              �?                                      @                                              @                                      �?       @       @       @                      �?      �?                                              �?                                      �?                                                      �?       @       @                                       @       @                                               @                                       @                                      �?                                       @      @      @                               @      @      �?                                      @      �?                                      @                                                      �?                               @       @                                       @      �?                                              �?                                       @                                                      �?                                                       @                                               @      �?      �?                                      �?      �?                                      �?                                                      �?                               @                �t�bub��+     hhubh)��}�(hhhhhNhKhKhG        hKhNhJQY%hG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKㅔh��B�1         �                    @���Ը��?�            `u@       [                     @ƒ_,���?�             n@       4       &             �?r��f?��?N            @^@       -                    �?&1��+��?*            @Q@                            �?��x�(��?             G@                           �?��S����?             ;@                           @9��8���?             8@              (             �?     ��?             0@	                           �?^N��)x�?             ,@
              '             �?9��8���?
             (@                           �?�8��8��?             @                            �?�q�q�?             @������������������������       �                      @������������������������       �                     �?              
             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?                           �?VUUUUU�?             @                           �?�Q����?             @                           @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @                           �?      �?              @                           �?�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     @!       (                    @6�80\��?             3@"       %                    �?��!pc�?             &@#       $                    �?�����H�?             "@������������������������       �                      @������������������������       �                     �?&       '                    �?      �?              @������������������������       �                     �?������������������������       �                     �?)       ,                     �?      �?              @*       +                    @z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @.       3                    @D%��N��?             7@/       0       
             �?X�<ݚ�?             "@������������������������       �                     @1       2                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     ,@5       R                    �?��]�`��?$             J@6       O                    �?�\��N��?             C@7       N       
             �?և���X�?             <@8       I                    �?
;&����?             7@9       H                    �?     ��?             0@:       E       "             �?��
ц��?
             *@;       >                    @���Q��?             $@<       =                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �??       D                     �?���Q��?             @@       A                    �?      �?             @������������������������       �                     �?B       C                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?F       G                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @J       M                    �?����X�?             @K       L                    �?r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @P       Q                    �?z�G�z�?             $@������������������������       �                      @������������������������       �                      @S       Z                    �?X�Cc�?
             ,@T       Y                    �?޾�z�<�?	             *@U       V       #             �?      �?             @������������������������       �                      @W       X                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@������������������������       �                     �?\       }                    @�7{`���?J            �]@]       h                    �?�����?#            �K@^       g                    �?
ףp=
�?             4@_       d                    �?F��ӭ��?             2@`       a       %             �?hE#߼�?             .@������������������������       �        	             &@b       c                    @      �?             @������������������������       �                     @������������������������       �                     �?e       f       !             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @i       z       %             �?���7F0�?            �A@j       u                    @@Q�f?��?             ?@k       r                    @ȵHPS!�?             :@l       m       "             �?���N8�?             5@������������������������       �                     0@n       q                    �?z�G�z�?             @o       p                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @s       t       )             �?���Q��?             @������������������������       �                     @������������������������       �                      @v       y                    �?{�G�z�?             @w       x                    @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @{       |                    @      �?             @������������������������       �                      @������������������������       �                      @~       �                    �?     0�?'             P@       �                    �?���GcT�?             C@�       �                    �?�m۶m��?             <@�       �       "             �?���ĳ��?	             .@�       �                    �?j�V���?             &@�       �       )             �?z�G�z�?             $@�       �       !             �?����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �       )             �?8�Z$���?             *@�       �                    �?      �?              @������������������������       �                     @�       �                    �?���Q��?             @�       �                    @      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    �?�z�G��?             $@������������������������       �                      @�       �                     @      �?              @�       �       &             �?      �?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �?��Q�}e�?             :@�       �                    @X��t��?             7@�       �       '             �?���7�?             6@�       �                    �?z�G�z�?             @������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        	             1@������������������������       �                     �?�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    @������?:            �Y@�       �                     @r�����?$            @P@�       �                    �?6?,R��?             B@�       �                    �?$I�$I��?             <@�       �                    �?�r����?             .@������������������������       �                     (@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                     �?�1G����?             *@������������������������       �                      @�       �                    @�x?r���?             &@�       �                    �?r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                    �?���Q��?             @������������������������       �                     @������������������������       �                      @�       �                    �?      �?              @������������������������       �                     �?�       �                    @����X�?             @������������������������       �                     @������������������������       �                      @�       �                    �?\B���?             =@�       �       &             �?r�q��?             8@�       �                    @�M�]��?             1@�       �       )             �?�����H�?             "@������������������������       �                     @�       �       	             �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                    �?����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                    �?����B�?            �B@�       �                    �?��f��?            �@@�       �                    �?\B���?             =@�       �                    �?H�7�&��?	             .@�       �       $             �?؇���X�?             ,@������������������������       �                     @�       �                    �?����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?�       �                     @T�r
^N�?	             ,@�       �                    @B{	�%��?             "@�       �                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�t�bh�h)h,K ��h.��R�(KK�KK��h�B�*       �C@     �I@      W@     �S@      M@      7@     �B@      I@      T@     �H@      1@      @      7@      6@      <@      >@      (@      @      @      @      2@      =@      (@      @      @      @      (@      *@      &@      @       @      @      @      "@      @      @       @      @      @      "@      @      @       @      @      @      @       @      @              @      @      @       @      @              @      @      �?       @      @                       @              �?      @                                      �?       @                                               @                                      �?                               @                      �?                       @                                                                      �?              @      �?      �?      �?                      @              �?      �?                      @              �?                              @                                                              �?                                                      �?                              �?                                                       @                       @                                                                      @       @                                      @       @                                               @                                      @                                               @                                                      @              �?              "@      @      @      �?      �?              "@      �?                                       @      �?                                       @                                                      �?                      �?              �?                              �?                                                              �?                                                      @      @      �?                                      @      �?                                              �?                                      @                                      @                                      @      0@      �?                              @       @      �?                              @                                                       @      �?                                       @                                                      �?                                      ,@                      4@      3@      $@      �?               @      4@      2@                                      (@      0@                                      (@      &@                                      @      "@                                      @      @                                      @      @                                      @      �?                                      @                                                      �?                                       @      @                                       @       @                                              �?                                       @      �?                                              �?                                       @                                                      �?                                      �?       @                                               @                                      �?                                                      @                                      @       @                                      @      �?                                              �?                                      @                                                      �?                                              @                                       @       @                                               @                                       @                                                      �?      $@      �?               @              �?      $@                       @              �?      �?                       @                                               @              �?      �?                                              �?                                      �?                                                      "@                                                      �?                      ,@      <@      J@      3@      @      �?      ,@      7@      "@      @      @      �?      &@              @               @      �?      &@              @               @      �?      &@              @                      �?      &@                                                              @                      �?                      @                                                                      �?                      �?               @                                               @                              �?                                               @                              @      7@      @      @       @              @      7@      �?       @       @              @      7@                                      �?      4@                                              0@                                      �?      @                                      �?      �?                                              �?                                      �?                                                      @                                       @      @                                              @                                       @                                                              �?       @       @                              �?               @                              �?                                                               @                                       @                                       @       @                                       @                                                       @                              @     �E@      .@      �?                      @      6@      *@                              @      3@      @                              �?       @      @                              �?       @       @                                       @       @                                      @       @                                      @                                                       @                                      @                                      �?                                                              @                               @      &@                                       @      @                                              @                                       @      @                                      �?      @                                      �?                                                      @                                      �?                                                      @                                              @      @                                               @                                      @      @                                      @      �?                                      �?      �?                                              �?                                      �?                                               @                                                      @                               @      5@       @      �?                              5@      �?      �?                              5@      �?                                      @      �?                                      @                                              �?      �?                                      �?                                                      �?                                      1@                                                              �?                       @              �?                               @                                                              �?                       @      �?      (@      >@     �D@      0@       @      �?      (@      9@      7@       @      �?      �?      $@      @      .@       @              �?      @      @      .@       @                                      *@       @                                      (@                                              �?       @                                      �?                                                       @              �?      @      @       @                                       @                              �?      @      @       @                      �?      @                                      �?                                                      @                                                      @       @                                      @                                                       @              �?              @       @                      �?                                                              @       @                                      @                                                       @                      �?               @      2@       @              �?               @      *@       @              �?                       @       @              �?                       @                                              @                      �?                      @                                              @                      �?                                                                               @                               @      @                                       @                                                      @                                              @                                              @      2@      ,@                              @      2@      $@                               @      1@      $@                              �?      (@       @                                      (@       @                                      @                                              @       @                                      @                                                       @                              �?                                              �?      @       @                              �?      �?      @                              �?      �?                                      �?                                                      �?                                                      @                                      @      �?                                              �?                                      @                                      @      �?                                              �?                                      @                                                              @�t�bubhhubh)��}�(hhhhhNhKhKhG        hKhNhJ��fbhG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK���h��B�#         ,                    �?.=T����?�            `u@              #             �?      �?3            �T@                           �?��R[s�?            �A@                           �?�>4և��?             <@                           �?ȵHPS!�?             :@������������������������       �        	             3@                           @և���X�?             @                           �?�q�q�?             @	                           �?z�G�z�?             @
                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                           @և���X�?             @                           �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @       #                    �?(���@��?            �G@                           �?�'�`d�?            �@@                            �?@4և���?
             ,@                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@       "       %             �?�����?
             3@              '             �?@4և���?             ,@������������������������       �                     $@        !                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @$       %       &             �?և���X�?	             ,@������������������������       �                      @&       +                     �?�q�q�?             (@'       (                    �?�q�q�?             @������������������������       �                     �?)       *                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @-       �                    @��� q�?�            @p@.       ]                    �?�:��X��?U            �a@/       L                    @p������?5            @U@0       K                    �?�	�FvD�?&             O@1       D                    �?�$I�$I�?#             L@2       ;       )             �?.�?�P��?             >@3       6                    �?����X�?	             ,@4       5                    �?ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@7       :                    �?      �?             @8       9                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @<       C                    �?     @�?             0@=       B                    �?X�Cc�?             ,@>       A                     @      �?              @?       @       
             �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                      @E       J                    �?$�q-�?             :@F       G                    �?`2U0*��?             9@������������������������       �                     6@H       I                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @M       \                    @P���� �?             7@N       S                     @>F?�!��?             5@O       P                    @      �?             @������������������������       �                      @Q       R       )             �?      �?              @������������������������       �                     �?������������������������       �                     �?T       [                    �?8߄*�u�?             1@U       V                    �?      �?
             0@������������������������       �                     *@W       Z                    �?�q�q�?             @X       Y                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @^       w       &             �?p����?              M@_       r                    �?�._�<�?            �B@`       o                    �?��ճC��?             6@a       j                    @�.�s�?             3@b       i       "             �?      �?             (@c       d                    �?"pc�
�?             &@������������������������       �                     @e       h                    �?�q�q�?             @f       g                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                     �?k       l                    �?����X�?             @������������������������       �                     @m       n                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @p       q       #             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @s       v                    @�.�?��?             .@t       u       "             �?r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@x       �                    @�a�a�?             5@y       �                    �?�$I�$I�?             @z       {                     �?{�G�z�?             @������������������������       �                     �?|                           @      �?             @}       ~                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     ,@�       �                    @�zq��?G            @]@�       �       
             �?�Ӫ�Ep�?             G@�       �                    @�%���^�?             2@�       �                    �?      �?
             (@�       �                    @      �?             @������������������������       �                      @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?      �?              @�       �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    @ �Cc}�?             <@������������������������       �                      @�       �                    �? ��WV�?             :@������������������������       �                     3@�       �                    �?؇���X�?             @������������������������       �                     @������������������������       �                     �?�       �                    @�,���=�?(            �Q@�       �       %             �?t��ճC�?             F@������������������������       �                     @������������������������       �                    �D@�       �                    �?�<ݚ�?             ;@������������������������       �                      @�       �                    �?�J�4�?             9@������������������������       �                     ,@�       �       $             �?���|���?             &@������������������������       �                     @������������������������       �                     @�t�bh�h)h,K ��h.��R�(KK�KK��h�B�        E@      G@     @S@      V@     �M@      >@     �D@     �D@                                      :@      "@                                      7@      @                                      7@      @                                      3@                                              @      @                                      @       @                                      @      �?                                       @      �?                                              �?                                       @                                               @                                                      �?                                              �?                                               @                                      @      @                                      �?      @                                              @                                      �?                                               @                                              .@      @@                                      @      :@                                      �?      *@                                      �?      �?                                              �?                                      �?                                                      (@                                      @      *@                                      �?      *@                                              $@                                      �?      @                                              @                                      �?                                              @                                               @      @                                               @                                       @      @                                       @      @                                      �?                                              �?      @                                              @                                      �?                                              @                                              �?      @     @S@      V@     �M@      >@      �?      @      Q@      I@      &@      "@                      E@     �B@      @                             �C@      5@       @                             �C@      .@       @                              .@      *@       @                              $@      @                                      "@      �?                                              �?                                      "@                                              �?      @                                      �?      �?                                      �?                                                      �?                                               @                                      @      "@       @                              @      "@                                      @      @                                      �?      @                                      �?                                                      @                                      @                                                      @                                                       @                              8@       @                                      8@      �?                                      6@                                               @      �?                                       @                                                      �?                                              �?                                              @                                      @      0@      @                              @      0@       @                               @      �?      �?                               @                                                      �?      �?                                      �?                                                      �?                              �?      .@      �?                                      .@      �?                                      *@                                               @      �?                                      �?      �?                                      �?                                                      �?                                      �?                                      �?                                                               @              �?      @      :@      *@      @      "@                      $@      *@      @      "@                      "@      @      @      @                      "@      @      @       @                      "@      @                                      "@       @                                      @                                              @       @                                       @       @                                               @                                       @                                               @                                                      �?                                                      @       @                                      @                                              �?       @                                      �?                                                       @                              �?               @                              �?                                                               @                      �?      "@              @                      �?                      @                      �?                                                                      @                              "@                      �?      @      0@                              �?      @       @                              �?       @       @                                      �?                                      �?      �?       @                              �?      �?                                      �?                                                      �?                                                       @                                       @                                                      ,@                                      �?      "@      C@      H@      5@              �?      "@     �A@      �?                      �?      @      $@      �?                      �?      @      @      �?                      �?       @              �?                               @                                      �?                      �?                      �?                                                                      �?                              @      @                                      �?      @                                              @                                      �?                                              @                                                      @                                      @      9@                                       @                                              �?      9@                                              3@                                      �?      @                                              @                                      �?                                                      @     �G@      5@                              @     �D@                                      @                                                     �D@                                              @      5@                                       @                                              @      5@                                              ,@                                      @      @                                              @                                      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hKhNhJ$�phG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKۅ�h��B�/         �                    �?��m4�?�            `u@       )                    �?Z$�����?�            @n@                           �?�ҿf���?1            �T@������������������������       �        
             (@       $                    �?\��_��?'            �Q@              $             �?Nd^����?"            �N@              
             �?8����?             G@                           �?`՟�G��?             ?@	                           �?��H�}�?             9@
                           �?��.k���?             1@                           �?      �?              @                           @      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @                           @�q�q�?             "@                            @      �?             @������������������������       �                      @              "             �?      �?             @������������������������       �                     �?                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @                           �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     .@       #                    �?������?	             .@       "                     �?�8��8��?             (@        !                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @%       &                    �?z�G�z�?             $@������������������������       �                     @'       (                    @      �?             @������������������������       �                      @������������������������       �                      @*       �                    �?>�����?f            �c@+       r                    �?��J���?H            �[@,       _                    @J:3�tK�?8            �U@-       V                    �?�J�)���?)            �O@.       E                    �?��8��x�?!             H@/       4                     �?��ׁsF�?             9@0       3                    �?VUUUUU�?             @1       2       !             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?5       8                    �? 9�����?             6@6       7                     @z�G�z�?             @������������������������       �                     �?������������������������       �                     @9       @                     @ҳ�wY;�?             1@:       ;       
             �?r�q��?
             (@������������������������       �                     @<       =       )             �?���Q��?             @������������������������       �                      @>       ?                    @�q�q�?             @������������������������       �                     �?������������������������       �                      @A       B       %             �?{�G�z�?             @������������������������       �                      @C       D                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?F       Q       "             �?l �&��?             7@G       L                    �?~h����?             ,@H       K                    �?�z�G��?             $@I       J                    �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @M       N                    �?      �?             @������������������������       �                     �?O       P       %             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?R       U                    �?X�<ݚ�?             "@S       T                    @����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @W       \       
             �?���Q��?             .@X       Y       %             �?$�q-�?             *@������������������������       �                     $@Z       [                     �?�q�q�?             @������������������������       �                     �?������������������������       �                      @]       ^                    �?      �?              @������������������������       �                     �?������������������������       �                     �?`       q       	             �?���x�?             7@a       n                    �?�z�G��?             4@b       e       %             �?،A��_�?             1@c       d                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @f       k                    @*x9/��?	             ,@g       j                    �?"pc�
�?             &@h       i                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @l       m                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?o       p                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @s       |       %             �?�q�q�?             8@t       u                    �?��(\���?             $@������������������������       �                     @v       {                    �?
ףp=
�?             @w       z                    �?VUUUUU�?             @x       y                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @}       ~                    �?؇���X�?	             ,@������������������������       �                     @       �                     @      �?              @�       �                    @؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �                    @�f��rL�?            �H@�       �                    �?�0OxJ'�?            �D@�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @�       �       (             �?N�y}IO�?            �B@�       �       &             �?�}�V`�?            �A@�       �                    �?
^N��)�?             <@�       �       #             �?���7�?             6@�       �                    @      �?              @�       �       )             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     ,@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     @�       �                    �?և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �                    �?      �?              @�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    @,��ݓ��?A             Y@�       �                    �?��?"m�?8             U@�       �       %             �?h��U�I�?,            �P@�       �                    �?l �&��?             7@�       �                     @      �?              @������������������������       �                      @������������������������       �                     @�       �       $             �?�Q����?
             .@�       �       
             �?ףp=
�?             $@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                     @���Q��?             @������������������������       �                      @������������������������       �                     @�       �                    @N��8��?            �E@�       �       !             �?���(\��?             $@�       �                    �?�$I�$I�?             @�       �       (             �?      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    @��Mu��?            �@@�       �                    @ȵHPS!�?             :@�       �                     �?���Q��?             @������������������������       �                      @������������������������       �                     @�       �                    @���N8�?             5@������������������������       �                     �?������������������������       �                     4@�       �                    �?և���X�?             @������������������������       �                     @������������������������       �                     @�       �                    �? )O��?             2@�       �                    @|	�%���?             "@������������������������       �                     @�       �                    �?VUUUUU�?             @������������������������       �                     �?�       �                     �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?X�<ݚ�?             "@�       �       %             �?؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                    �?     ��?	             0@�       �                    �?VUUUUU�?             "@�       �                    �?�Q����?             @������������������������       �                     �?�       �                    �?      �?             @������������������������       �                      @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�t�bh�h)h,K ��h.��R�(KK�KK��h�B)        I@     �L@     �Q@     �T@     �J@      =@      G@      F@      I@     �N@      9@      0@     �F@      C@                                      (@                                             �@@      C@                                      9@      B@                                      ,@      @@                                      ,@      1@                                      "@      0@                                      "@       @                                      @       @                                       @       @                                               @                                       @                                              @                                              @      @                                      @      @                                               @                                      @      �?                                      �?                                               @      �?                                              �?                                       @                                                      @                                               @                                      @      �?                                      @                                                      �?                                              .@                                      &@      @                                      &@      �?                                      @      �?                                      @                                                      �?                                      @                                                      @                                       @       @                                      @                                               @       @                                               @                                       @                                              �?      @      I@     �N@      9@      0@      �?      @      D@     �@@      1@      ,@              @     �A@      3@      1@      &@               @     �@@      .@       @      @              �?      4@      ,@       @      @              �?      *@      @      @      �?              �?                      �?      �?              �?                      �?                                              �?                      �?                                                                              �?                      *@      @      @                              �?              @                              �?                                                              @                              (@      @       @                              $@       @                                      @                                              @       @                                       @                                              �?       @                                      �?                                                       @                                       @      �?       @                               @                                                      �?       @                                               @                                      �?                                      @      &@      �?      @                      @      @      �?                              @      @                                       @      @                                       @                                                      @                                      @                                                      @      �?                                      �?                                               @      �?                                       @                                                      �?                                      @              @                              @               @                              @                                                               @                                               @              �?      *@      �?                              �?      (@                                              $@                                      �?       @                                      �?                                                       @                                              �?      �?                                              �?                                      �?                                       @       @      @      "@      @               @       @      @      "@      @               @              @      "@       @               @              �?                                              �?                               @                                                              @      "@       @                               @      "@                                       @      �?                                       @                                                      �?                                               @                                      �?               @                                               @                              �?                                       @                      �?                       @                                                                      �?                                              @      �?      �?      @      ,@              @      �?      �?      @       @              �?                      @                              �?      �?               @              �?      �?      �?                              �?      �?                                      �?      �?                                                                                      �?              �?                                                               @                                              (@               @                              @                                              @               @                              @              �?                              @                                                              �?                                              �?              �?      $@      <@       @       @              �?      $@      <@       @                               @               @                                               @                               @                                      �?       @      <@                              �?      @      <@                              �?      @      8@                              �?              5@                              �?              @                              �?               @                              �?                                                               @                                              @                                              ,@                                      @      @                                      @                                                      @                                      @      @                                      @                                                      @                                       @                                                              @       @                                       @       @                                       @                                                       @                                      @              @      *@      4@      6@      <@      *@              (@      4@      3@      ;@      @              @      *@      1@      :@      @              @      "@      "@                               @              @                               @                                                              @                              @      "@      @                              �?      "@                                      �?      @                                              @                                      �?                                                      @                                       @              @                               @                                                              @                              �?      @       @      :@      @              �?      @      @                              �?      @       @                              �?      @                                              @                                      �?                                                      �?       @                                      �?                                                       @                                              @                                              @      :@      @                              @      7@                                       @      @                                       @                                                      @                                      �?      4@                                      �?                                                      4@                                              @      @                                              @                                      @                      @      @       @      �?       @              @      �?      �?      �?                      @                                                      �?      �?      �?                                      �?                                      �?              �?                                              �?                              �?                                              @      �?               @                      @      �?                                      @                                                      �?                                                               @      @      �?              @      �?      @      @      �?              @      �?                      �?              @      �?                      �?                                                              @      �?                                       @                                              �?      �?                                      �?                                                      �?              @                                                                                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hKhNhJW:+LhG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKم�h��Bx/         t       &             �?������?�            `u@       K                    �?O�
@�?v            �g@       $       
             �?�?�P�a�?N             ^@                           �?     ��?&             P@       
                    �?���.�?
             3@       	                    �?      �?             0@              (             �?��S�ۿ?             .@������������������������       �                     ,@������������������������       �                     �?������������������������       �                     �?                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?                           �?t�����?            �F@                           @�p9W���?
             3@������������������������       �                     @                           @pƵHP�?             *@������������������������       �                     @                           @      �?             @������������������������       �                     @������������������������       �                     @                           �?h��9J�?             :@                           @��ˠ�?             &@������������������������       �                     @                           �?������?             @������������������������       �                     @                           �?      �?             @������������������������       �                     @������������������������       �                     �?       #                    @ƒ_,���?             .@       "                    �?z�G�z�?             $@        !                    @�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @%       >                    �?4և����?(             L@&       =                     @0�@g���?            �D@'       (                    �?��[��"�?             B@������������������������       �                      @)       .                    �?k��\��?             A@*       +                    �?"pc�
�?             &@������������������������       �                      @,       -                    @�q�q�?             @������������������������       �                     �?������������������������       �                      @/       6                    @�\@˜��?             7@0       5                     @���Q��?             .@1       4                    �?      �?             (@2       3                    @���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @7       <                    @      �?              @8       9                    �?�q�q�?             @������������������������       �                     @:       ;                    @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @?       @                    @ƒ_,���?	             .@������������������������       �                      @A       D                    �?�n_Y�K�?             *@B       C                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @E       J                    �?      �?              @F       I                    �?      �?             @G       H                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @L       o       (             �?�/â���?(            @Q@M       ^       '             �?Z.ҫ; �?%             O@N       S                    @1�rXQ�?            �B@O       R                      @��Q��?             $@P       Q                    @և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @T       Y                    @a�J�GT�?             ;@U       X                    �?z�G�z�?             @V       W                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @Z       ]       "             �?�eP*L��?             6@[       \                    @p�ݯ��?             3@������������������������       �                     (@������������������������       �                     @������������������������       �                     @_       n                    �?46<��?             9@`       k                    �?x�5?,R�?             2@a       j                    �?*D>��?	             *@b       g                    @��(\���?             $@c       d       #             �?      �?              @������������������������       �                     @e       f                    �?      �?             @������������������������       �                     @������������������������       �                     �?h       i                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @l       m                     @���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @p       s                    �?�$I�$I�?             @q       r                    @z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @u       �                    �?8]��"�?j             c@v       �                    �?��j�9��?Z            @`@w       �                    @Ӆ��?L            �Z@x                           �?2����}�?%            �F@y       z                    �?X�Cc�?             ,@������������������������       �                      @{       |                    @�������?
             (@������������������������       �                     $@}       ~                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @@�sP�?             ?@�       �                    �?x?r����?             6@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?ףp=
�?             4@������������������������       �                     &@�       �                    �?�<ݚ�?	             "@������������������������       �                      @�       �                    �?����X�?             @�       �                    �?      �?             @�       �                     @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �?��E���?             "@�       �                     @�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                     �?r�q��?             @�       �                    �?      �?             @������������������������       �                      @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    �?v��V:e�?'             O@�       �       
             �?���Q��?             $@������������������������       �                     @������������������������       �                     @�       �                    @n_Y�K�?!             J@�       �                    �?�$c���?            �D@������������������������       �                     �?�       �                    �?z�G�z�?             D@�       �                    �?$�q-�?             :@������������������������       �                     7@�       �                     @�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �       "             �?X�Cc�?             ,@�       �       '             �?"pc�
�?             &@������������������������       �                     @�       �                    @      �?              @�       �                    �?      �?             @�       �       !             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                    @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    @������?             &@�       �                    �?      �?              @�       �                    �?r�q��?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �?8��Moz�?             7@������������������������       �                     @�       �                    �?tk~X��?             2@������������������������       �        	             *@�       �       '             �?���Q��?             @������������������������       �                     @������������������������       �                      @�       �                    �?��;5r�?             7@�       �                    �?      �?              @�       �                    �?r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @ƒ_,���?             .@������������������������       �                     @�       �                    @ףp=
��?             $@�       �                    �?      �?             @������������������������       �                     �?�       �                    @�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?�t�b�x     h�h)h,K ��h.��R�(KK�KK��h�B�(        ?@     �J@     �U@     �V@     �G@      A@      @      @      E@     �O@     �F@      =@       @      @     �A@      F@      8@      &@       @      @      =@      3@       @       @              �?      .@      �?               @              �?      ,@      �?                                      ,@      �?                                      ,@                                                      �?                              �?                                                      �?                       @                                               @                      �?                               @      @      ,@      2@       @                              "@      @      @                              @                                              @      @      @                                      @                                      @              @                                              @                              @                               @      @      @      &@      @                      @      @      @                                      @                                      @      �?      @                              @                                                      �?      @                                              @                                      �?                               @                       @      @               @                       @                      �?                       @                                               @                      �?                                              �?                                                                              @                              @      9@      0@      "@                      @      7@       @      @                      @      2@       @      @                                       @                              @      2@      @      @                              "@       @                                       @                                              �?       @                                      �?                                                       @                              @      "@      @      @                      @      "@                                      @      "@                                      @       @                                      @                                                       @                                              @                                      @                                                              @      @                                       @      @                                              @                                       @      �?                                              �?                                       @                                               @                                      @                                               @       @      @                               @                                                       @      @                                      �?      @                                      �?                                                      @                                      @      �?                                      @      �?                                      �?      �?                                      �?                                                      �?                                       @                                              @              @              @      3@      5@      2@                      @      3@      4@      0@                      @      @      0@      *@                      @      @              @                      @                      @                      @                                                                      @                              @                                              �?      0@      $@                              �?      @                                      �?      �?                                      �?                                                      �?                                              @                                              (@      $@                                      (@      @                                      (@                                                      @                                              @                      @      .@      @      @                      @       @      @      @                      �?       @      �?      @                      �?       @      �?                              �?      @                                              @                                      �?      @                                              @                                      �?                                                      �?      �?                                              �?                                      �?                                                              @                       @              @                               @                                                              @                                      @                      @                              �?       @      @                              �?              @                                                                              �?                                                       @      9@     �H@     �F@      ;@       @      @      6@      D@      F@      1@       @      @      1@      ;@     �D@      .@       @      @      *@      5@      @       @      �?      �?      $@       @      �?                      �?               @                                      $@              �?                      �?      $@                                                              �?                      �?                      �?                                                                      �?      @      3@      @       @      �?              @      2@      �?                              �?              �?                                              �?                              �?                                               @      2@                                              &@                                       @      @                                               @                                       @      @                                       @       @                                       @      �?                                              �?                                       @                                                      �?                                              @                                              �?      @       @      �?                      �?               @                              �?                                                               @                                      @              �?                              @              �?                               @                                              �?              �?                                              �?                              �?                                               @                              @      @      A@      *@      �?      @      @      @                                              @                                      @                                                              A@      *@      �?      @                     �@@      @              �?                                              �?                     �@@      @                                      8@       @                                      7@                                              �?       @                                      �?                                                       @                                      "@      @                                      "@       @                                      @                                              @       @                                      @      �?                                       @      �?                                       @                                                      �?                                      �?                                              @      �?                                      @                                                      �?                                              @                                      �?      @      �?      @                      �?      @      �?                              �?      @                                      �?      �?                                      �?                                                      �?                                              @                                              �?      �?                                      �?                                                      �?                                                      @      @      *@      @       @                      @                                                      *@      @       @                              *@                                                      @       @                                      @                                                       @                      @      "@      �?      $@                      �?      �?      �?      @                      �?                      @                      �?                                                                      @                              �?      �?                                      �?                                                      �?                               @       @              @                              @                                       @      @              @                       @       @                                              �?                                       @      �?                                              �?                                       @                                                      �?              @                                              @                              �?                                �t�bubhhubh)��}�(hhhhhNhKhKhG        hKhNhJF<KdhG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKυ�h��BH-         2                    �?�"�|��?�            `u@                           �?7�A�0�?<             V@������������������������       �                     1@       -                    �?��M��?1            �Q@                            �?�θ�?,            @P@                           @�iʫ{�?"            �J@                           �?�KM�]�?             C@              !             �?�J�4�?             9@	              "             �?d}h���?             ,@
                           �?�C��2(�?	             &@������������������������       �                      @              	             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?                           �?�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@������������������������       �                     *@              %             �?�q�q�?             .@                           �?r�q��?             (@������������������������       �                     @              )             �?����X�?             @                           @z�G�z�?             @������������������������       �                     @������������������������       �                     �?              "             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @!       ,                    �?      �?
             (@"       %       )             �?���Q��?             $@#       $       &             �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @&       +       $             �?���Q��?             @'       (       
             �?      �?             @������������������������       �                      @)       *                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @.       1                     �?r�q��?             @/       0                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @3       �       
             �?&���*�?�            �o@4       �                    �?4�$q��?R            �`@5       n                    �?y���?I            �]@6       I       %             �?��1M�?+            @P@7       B                    �?�2�tk~�?             2@8       A                    �?      �?              @9       @                    �?VUUUUU�?             @:       =                    @      �?             @;       <                    �?      �?              @������������������������       �                     �?������������������������       �                     �?>       ?       "             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @C       H                    �?ףp=
��?             $@D       G       )             �?�8��8��?             @E       F                     @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @J       W                    �?T�#�3@�?            �G@K       V                    �?��2Tv�?
             .@L       S                    �?�θ�?	             *@M       R                    �?ףp=
��?             $@N       O                    @x�5?,�?             "@������������������������       �                     @P       Q                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?T       U       (             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @X       e                    �?     @�?             @@Y       b       	             �?x��J��?             7@Z       ]                    �?�a�a�?             5@[       \                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?^       _                    �?�����H�?	             2@������������������������       �                     &@`       a                    �?����X�?             @������������������������       �                     @������������������������       �                      @c       d                    @      �?              @������������������������       �                     �?������������������������       �                     �?f       m       "             �?��"e���?             "@g       h                    @������?             @������������������������       �                     �?i       j       	             �?      �?             @������������������������       �                      @k       l                    @      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @o       x                    �?�8�l��?            �J@p       u                    @��!pc�?            �@@q       t                     �?�%d���?             =@r       s                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     ;@v       w       &             �?      �?             @������������������������       �                     @������������������������       �                     �?y       |                    �?p=
ףp�?             4@z       {                    @z�G�z�?             @������������������������       �                     @������������������������       �                     �?}       �       )             �?�q�q�?             .@~              &             �?�eP*L��?             &@������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    @�r����?	             .@������������������������       �                     (@�       �       '             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    @�=��R�?N            @^@�       �                     @ū\��5�?.            �P@�       �                    �?ĨS@Q��?)            �N@�       �                    �?6M5���?            �D@�       �                    �?޾�z�<�?             *@�       �                    �?�$I�$I�?             @�       �                    �?      �?             @������������������������       �                     �?�       �       $             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                    @և���X�?             <@������������������������       �                     "@�       �                    �?p�ݯ��?             3@�       �                    �?d}h���?             ,@������������������������       �                      @�       �       '             �?      �?             @������������������������       �                      @�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    �?H�z�G�?             4@������������������������       �                     �?�       �                    @�d�����?             3@������������������������       �                     �?�       �       	             �?�X�<ݺ?             2@������������������������       �        
             1@������������������������       �                     �?�       �                    �?�q�q�?             @�       �       #             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �       &             �?��h]���?              K@�       �                    �?TR'����?             I@�       �                    �?9��8�#�?             H@�       �                     @�E��ӭ�?
             2@�       �                    �?$�q-�?             *@������������������������       �                     @�       �       '             �?؇���X�?             @������������������������       �                     �?������������������������       �                     @�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                    �?H�z�G�?             >@�       �                    �?V��6���?             1@������������������������       �                     �?�       �                    �?     ��?             0@�       �                    �?�����H�?             "@������������������������       �                      @������������������������       �                     �?�       �                    @����X�?             @�       �       $             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �?�	j*D�?             *@�       �                    �?���Q��?             $@�       �                    �?�q�q�?             @�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     @�t�bh�h)h,K ��h.��R�(KK�KK��h�B�&        C@     �N@     @U@     @V@      F@      9@     �B@     �I@                                      1@                                              4@     �I@                                      .@      I@                                      "@      F@                                      @      A@                                      @      5@                                      @      &@                                      �?      $@                                               @                                      �?       @                                      �?                                                       @                                       @      �?                                       @                                                      �?                                      �?      $@                                      �?                                                      $@                                              *@                                      @      $@                                       @      $@                                              @                                       @      @                                      �?      @                                              @                                      �?                                              �?      �?                                              �?                                      �?                                              @                                              @      @                                      @      @                                      @      �?                                              �?                                      @                                               @      @                                      �?      @                                               @                                      �?      �?                                      �?                                                      �?                                      �?                                                       @                                      @      �?                                      @      �?                                              �?                                      @                                               @                                              �?      $@     @U@     @V@      F@      9@      �?      "@      O@     �B@      (@      (@      �?      "@     �H@     �A@      (@      (@      �?      @      *@      9@      &@      &@      �?       @      @      @      �?      @      �?              �?              �?      @      �?              �?              �?      @      �?              �?              �?      �?      �?              �?                                              �?                              �?                                                                              �?      �?                                      �?                                                      �?                                               @                                               @               @      @      @                               @      �?      @                               @      �?                                       @                                                      �?                                                      @                                      @                                       @      @      6@      $@      @               @      @      @       @       @               @      @      @               @                      @      @               @                      @      @              �?                      @                                                      @              �?                                              �?                              @                                                              �?               @              �?                               @                                                              �?                                                       @                               @      2@       @      @                      �?      0@      @      �?                      �?      0@      @                              �?               @                                               @                              �?                                                      0@       @                                      &@                                              @       @                                      @                                                       @                                              �?      �?                                      �?                                                      �?                      �?       @      @      @                      �?              @      @                      �?                                                              @      @                                       @                                              �?      @                                      �?                                                      @                               @                              @      B@      $@      �?      �?              @      ;@              �?      �?              �?      ;@                      �?              �?                              �?              �?                                                                              �?                      ;@                                      @                      �?                      @                                                                      �?                      �?      "@      $@                              �?      @                                              @                                      �?                                                      @      $@                                      @      @                                              @                                      @                                                      @                                      *@       @                                      (@                                              �?       @                                      �?                                                       @                              �?      7@      J@      @@      *@              �?      7@     �D@       @                      �?      3@     �C@       @                              2@      6@      �?                               @      $@      �?                               @      @      �?                               @      �?      �?                                      �?                                       @              �?                                              �?                               @                                                      @                                              @                                      0@      (@                                      "@                                              @      (@                                      @      &@                                               @                                      @      @                                               @                                      @      �?                                              �?                                      @                                              @      �?                                      @                                                      �?                              �?      �?      1@      �?                                              �?                      �?      �?      1@                              �?                                                      �?      1@                                              1@                                      �?                                              @       @                                      �?       @                                      �?                                                       @                                      @                                                      &@      >@      *@                              @      >@      *@                              @      >@      &@                              @      *@                                      �?      (@                                              @                                      �?      @                                      �?                                                      @                                      @      �?                                              �?                                      @                                               @      1@      &@                               @      *@       @                                              �?                               @      *@      �?                                       @      �?                                       @                                                      �?                               @      @                                       @      �?                                       @                                                      �?                                              @                                              @      "@                                      @      @                                      @       @                                       @       @                                       @                                                       @                                       @                                                      @                                              @                                               @                              @                �t�bubhhubh)��}�(hhhhhNhKhKhG        hKhNhJؽ�hG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK���h��Bh%         T       %             �?�ƄҢ*�?�            `u@       	                    �?lb	�?c             c@                           @�?             1@������������������������       �        	             (@                           �?{�G�z�?             @������������������������       �                      @                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @
       C       
             �?jiiiii�?W             a@       2                    �?�L�p�?6             U@       #       !             �?2Y�Qo��?!             K@                            @��&����?            �B@                           �?��[r��?             5@                           �?���Q��?             .@                           �?ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@                           �?z�G�z�?             @������������������������       �                      @                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @                           �?r�q��?             @������������������������       �                     �?������������������������       �                     @       "                    �?     @�?             0@                           �?>;n,��?             &@������������������������       �                     @       !                    @0�����?             @                            �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @$       +                    @k��\��?
             1@%       &                    �?j�V���?             &@������������������������       �                      @'       *                    �?�����H�?             "@(       )                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @,       -                    �?      �?             @������������������������       �                     �?.       1                    �?z�G�z�?             @/       0                     @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @3       <                    �?�h$���?             >@4       ;                    �?��S���?
             .@5       6                    �?�q�q�?             (@������������������������       �                     @7       :                    �?����X�?             @8       9                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @=       >                    �?�.�?��?             .@������������������������       �                     @?       B                     �?��!pc�?             &@@       A                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@D       S                    @��WV��?!             J@E       N                    �?X1��^�?             E@F       I                    @b�2�tk�?             2@G       H                    �?      �?             (@������������������������       �                     "@������������������������       �                     @J       M                    �?�q�q�?             @K       L       $             �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?O       P                    @r�q��?             8@������������������������       �                     0@Q       R                    �?      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     $@U       �                    @FR���?s            �g@V       y                    �?�2��,��?5            �V@W       p                    �?���Y��?,            �S@X       o                    @�'N��?#            �N@Y       h                    �?H�z�G�?             D@Z       c                    �?���>4��?             <@[       b                    �?���|���?             6@\       a                    �?և���X�?             ,@]       ^       #             �?      �?
             (@������������������������       �                     @_       `                    �?؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                      @d       e       '             �?r�q��?             @������������������������       �                     @f       g                    �?      �?              @������������������������       �                     �?������������������������       �                     �?i       j                     @r�q��?             (@������������������������       �                     �?k       n                    �?�C��2(�?             &@l       m                      @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@������������������������       �                     5@q       x                    �?P�|�@�?	             1@r       s       '             �?�1G����?             *@������������������������       �                     @t       u                    �?      �?              @������������������������       �                     @v       w                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @z       {                    �?;�;��?	             *@������������������������       �                     @|       }                    �?      �?              @������������������������       �                     @~                           �?      �?             @������������������������       �                     �?�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    @jw�3=�?>            �X@�       �                    �?�T`�[k�?%            �J@�       �                    @8��8���?"             H@�       �                    �?�q�q�?             8@�       �                    @���Q��?
             .@�       �                    �?      �?              @������������������������       �                     �?�       �                    �?؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �       $             �?�����H�?             "@�       �                    �?      �?             @������������������������       �                      @�       �       )             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     8@������������������������       �                     @�       �                    �?f.i��n�?            �F@�       �       )             �?`՟�G��?             ?@�       �                    �?�t����?	             1@�       �                    �?      �?             0@�       �                    �?z�G�z�?             .@�       �                    @؇���X�?             ,@������������������������       �                     &@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                    �?؇���X�?             ,@�       �                    �?�q�q�?             @�       �                     �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                     ,@�t�bh�h)h,K ��h.��R�(KK�KK��h�B         E@     �J@     �Q@     �U@      M@     �@@     �A@      H@      E@      7@      @       @      (@               @               @      �?      (@                                                               @               @      �?                                       @                               @                      �?                                              �?                       @                              7@      H@      D@      7@      �?      �?      0@     �B@      4@      "@      �?      �?      "@      <@      &@      @      �?      �?      @      3@      &@                               @      "@      $@                              �?      @      $@                              �?              "@                              �?                                                              "@                                      @      �?                                       @                                               @      �?                                              �?                                       @                                      �?      @                                      �?                                                      @                                      @      $@      �?                              @      @      �?                                      @                                      @      �?      �?                              @      �?                                      @                                                      �?                                                      �?                                      @                                       @      "@              @      �?      �?       @       @                      �?               @                                                       @                      �?                      @                      �?                      @                                                                      �?                      @                                              �?              @              �?              �?                                                              @              �?                               @              �?                               @                                                              �?                               @                      @      "@      "@      @                      @       @                                      @      @                                      @                                               @      @                                       @      �?                                       @                                                      �?                                              @                                              @                                              �?      "@      @                                              @                              �?      "@      �?                              �?              �?                              �?                                                              �?                                      "@                              @      &@      4@      ,@                      @      &@      4@      @                      @      &@                                      @      "@                                              "@                                      @                                              @       @                                      @      �?                                              �?                                      @                                                      �?                                                      4@      @                                      0@                                              @      @                                              @                                      @                                                      $@                      @      @      <@     �O@     �K@      ?@      @      @      <@     �I@                       @      @      6@     �H@                                      1@      F@                                      1@      7@                                      .@      *@                                      ,@       @                                      @       @                                      @      @                                              @                                      @      �?                                      @                                                      �?                                               @                                       @                                              �?      @                                              @                                      �?      �?                                      �?                                                      �?                                       @      $@                                      �?                                              �?      $@                                      �?      �?                                      �?                                                      �?                                              "@                                              5@                       @      @      @      @                       @      �?      @      @                                              @                       @      �?      @                                              @                               @      �?                                              �?                                       @                                                      @                                      @              @       @                      @                                                              @       @                                      @                                               @       @                                      �?                                              �?       @                                      �?                                                       @                                              (@     �K@      ?@                              (@     �D@                                      @     �D@                                      @      1@                                      @      "@                                      @       @                                              �?                                      @      �?                                              �?                                      @                                                      @                                      �?       @                                      �?      @                                               @                                      �?      �?                                              �?                                      �?                                                      @                                              8@                                      @                                                      ,@      ?@                                      ,@      1@                                      (@      @                                      (@      @                                      (@      @                                      (@       @                                      &@                                              �?       @                                      �?                                                       @                                              �?                                              �?                                              �?                                       @      (@                                       @      @                                       @       @                                               @                                       @                                                       @                                               @                                              ,@�t�bubhhubh)��}�(hhhhhNhKhKhG        hKhNhJX��vhG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKم�h��Bx/         �                    @�a'��?�            `u@       Y                    �?\!�ab�?�            �k@       >                    @6��?�)�?P            �`@              %             �?���V�/�?9             Y@                           �?V"H�~�?            �E@                           �?���Q��?             D@       
                    @     0�?             @@       	                    �?d}h���?
             ,@������������������������       �                     @������������������������       �        	             &@                           �?0�����?	             2@������������������������       �                     �?                           �?�IєX�?             1@������������������������       �                     (@              
             �?z�G�z�?             @              )             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @                           �?      �?              @������������������������       �                     �?                           �?և���X�?             @������������������������       �                      @              $             �?���Q��?             @������������������������       �                     @������������������������       �                      @                           @�q�q�?             @������������������������       �                     �?                           �?      �?              @������������������������       �                     �?������������������������       �                     �?        -                    @��y��?            �L@!       ,       )             �?�q�q�?             8@"       %                    �?ҳ�wY;�?
             1@#       $                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?&       )                    �?����S�?             ,@'       (       	             �?�8��8��?             (@������������������������       �                     &@������������������������       �                     �?*       +                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @.       7                    �?8�#�(�?            �@@/       4                    �?ҳ�wY;�?             1@0       3                    �?޾�z�<�?             *@1       2                    �?r�q��?             (@������������������������       �                     $@������������������������       �                      @������������������������       �                     �?5       6       '             �?      �?             @������������������������       �                      @������������������������       �                      @8       =                    �?     ��?             0@9       <                     �?�$I�$I�?             @:       ;                     @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     "@?       L                    �?6c����?             A@@       K                    �?r�q��?	             (@A       H       %             �?4և����?             @B       E                    �?      �?             @C       D                    �?      �?              @������������������������       �                     �?������������������������       �                     �?F       G       $             �?      �?              @������������������������       �                     �?������������������������       �                     �?I       J                     @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @M       X                    �?��eP*L�?             6@N       S                    �?b>���?             5@O       P                    �?�r����?	             .@������������������������       �                     �?Q       R                    @@4և���?             ,@������������������������       �                     *@������������������������       �                     �?T       W                    �?�8��8��?             @U       V       
             �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?Z       i                    �?����?8            @V@[       \                    �?���@M^�?             ?@������������������������       �        	             ,@]       ^                    �?�t����?
             1@������������������������       �                      @_       h                    �?z�G�z�?	             .@`       a                     �?���!pc�?             &@������������������������       �                     @b       g                    �?և���X�?             @c       d       #             �?      �?             @������������������������       �                      @e       f                     @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @j       �       
             �?~Riv���?%             M@k       x                    �?ףp=
��?             D@l       s       "             �?v�f��?             1@m       r       )             �?x�5?,�?             "@n       o                    �?�8��8��?             @������������������������       �                      @p       q                    @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @t       u                    �?      �?              @������������������������       �                     @v       w                     �?�q�q�?             @������������������������       �                     �?������������������������       �                      @y       �       %             �?x��J��?             7@z       �                    @.y0��k�?
             *@{       �       )             �?�8��8��?	             (@|       }                    �?؇���X�?             @������������������������       �                     @~                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                    �?      �?             $@������������������������       �                     @�       �                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    �?�8��8��?
             2@�       �                    �?���Q��?             .@�       �                    �?޾�z�<�?             *@�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @�       �       )             �?�����H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    �?�
�OK��?K            �]@�       �       &             �?�q�q,�?>             X@�       �                    @8�&���?'             N@�       �                    �?���^�?             ;@�       �                    �?�KM�]�?             3@�       �                    @      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     .@�       �                    �?      �?              @������������������������       �                     @������������������������       �                     @�       �                    @6YE�?            �@@�       �                    �?ȵHPS!�?             :@������������������������       �                     7@������������������������       �                     @�       �                    �?����X�?             @������������������������       �                      @������������������������       �                     @�       �       )             �?uk~X��?             B@�       �                     @UUUUUU�?             (@�       �                    @�q�q�?             @�       �       (             �?      �?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �       #             �?      �?             @������������������������       �                     �?�       �       
             �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                     �?r�q��?             8@�       �       $             �?@�0�!��?	             1@�       �                    �?�q�q�?             (@������������������������       �                     �?�       �                    @���!pc�?             &@�       �                    �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                    �?{�G�z�?             @������������������������       �                      @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?�$I�$I�?             @�       �                    �?{�G�z�?             @�       �                    @      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                    �?p�u=q��?             7@�       �       !             �?
ц�s�?             *@�       �                    @�<ݚ�?             "@������������������������       �                     @�       �       %             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @�       �       &             �?���(\��?             $@�       �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @�t�bh�h)h,K ��h.��R�(KK�KK��h�B�(       �G@      J@      T@      U@     �N@      2@      :@      A@     �P@      K@      >@      (@      @      2@      F@     �C@      8@      @      @      0@      E@      6@      .@              @      ,@      3@      @                      @      *@      3@      @                      @      (@      0@      �?                      @      &@                                      @                                                      &@                                              �?      0@      �?                              �?                                                      0@      �?                                      (@                                              @      �?                                       @      �?                                       @                                                      �?                                       @                                      �?      @      @                              �?                                                      @      @                                               @                                      @       @                                      @                                                       @                       @      �?                                      �?                                              �?      �?                                      �?                                                      �?                                               @      7@      1@      .@                       @      3@      @                               @      (@      @                              �?               @                                               @                              �?                                              �?      (@      �?                                      &@      �?                                      &@                                                      �?                              �?      �?                                              �?                                      �?                                                      @                                              @      ,@      .@                              @      (@       @                              �?      $@       @                                      $@       @                                      $@                                                       @                              �?                                               @       @                                       @                                                       @                                      �?       @      *@                              �?       @      @                              �?       @                                      �?                                                       @                                                      @                                              "@                       @       @      1@      "@      @              �?       @      �?      @       @              �?       @      �?      �?       @              �?       @      �?                                      �?      �?                                      �?                                                      �?                              �?      �?                                              �?                                      �?                                                                      �?       @                                               @                                      �?                                              @                      �?              0@      @       @              �?              0@       @       @                              *@       @                                              �?                                      *@      �?                                      *@                                                      �?                      �?              @               @                              @               @                              @                                                               @              �?                                                                      �?              5@      0@      7@      .@      @       @      3@      (@                                      ,@                                              @      (@                                       @                                              @      (@                                      @       @                                              @                                      @      @                                      @      �?                                       @                                              �?      �?                                              �?                                      �?                                                      @                                              @                                       @      @      7@      .@      @       @       @      @      6@      @       @      @       @      @      @              �?      @              @      @              �?                      @       @              �?                               @                                      @                      �?                      @                                                                      �?                              @                               @              �?                      @                                              @       @              �?                                              �?                               @                                                      �?      0@      @      �?                      �?      &@              �?                      �?      &@                                      �?      @                                              @                                      �?       @                                      �?                                                       @                                              @                                                              �?                              @      @                                              @                                      @      �?                                      @                                                      �?                                      �?      $@      @      @                      �?      $@      @                              �?      $@       @                                       @       @                                               @                                       @                                      �?       @                                      �?                                                       @                                                       @                                                      @      5@      2@      *@      >@      ?@      @      ,@      $@      &@      <@      ;@      @       @              @      9@      9@      @       @              @      6@                       @                      1@                       @                       @                       @                                                                       @                                              .@                                      @      @                                      @                                                      @                                              @      9@      @                              @      7@                                              7@                                      @                                                       @      @                                       @                                                      @      (@      $@       @      @       @      �?      �?       @      @       @       @      �?      �?       @              �?       @              �?       @              �?                      �?                      �?                                              �?                      �?                                                       @                                                                       @                              @      �?              �?                              �?                                      @                      �?                                              �?                      @                              &@       @      @      �?                      $@      @       @      �?                       @      @                                              �?                                       @      @                                       @      @                                              @                                       @                                              @                                               @               @      �?                                       @                               @                      �?                       @                                                                      �?                      �?      @       @                              �?       @       @                                       @       @                                               @                                       @                                      �?                                                       @                                      @       @       @       @      @               @      @       @       @                              @               @                              @                                              �?               @                              �?                                                               @                       @               @                                               @                               @                                              @      �?                      @              �?                              @                                              @              �?                                              @      �?                                              �?                                      @                                        �t�bub�?     hhubh)��}�(hhhhhNhKhKhG        hKhNhJ���EhG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKۅ�h��B�/         j       %             �?�`�����?�            `u@                           �?���:��?`            @c@                           �?�n����?
             2@                           �?�θ�?             *@                           �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@	       
                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @       7                    �?�V�e�t�?V             a@       "       '             �?     |�?'             P@                           �?z�;c��?             =@              
             �?��1G���?             :@                           �?Y�����?             &@                            �?X�<ݚ�?             "@                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?                           �?r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @                           @�Q����?             .@                           �?      �?             @������������������������       �                      @                           �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     "@        !                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?#       (                    @�~VDq�?            �A@$       '                    �?�q�q�?             @%       &                    �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?)       2                     �?$:9$A��?             =@*       +                    �?8��8���?             8@������������������������       �                     *@,       /       
             �?j�V���?             &@-       .                    �?      �?              @������������������������       �                     �?������������������������       �                     �?0       1                    �?�����H�?             "@������������������������       �                     �?������������������������       �                      @3       6                    �?���Q��?             @4       5                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?8       _                    �?n�����?/             R@9       Z                    �?6д>���?%             M@:       O                    �?E3����?"             K@;       H                    �?_j����?             C@<       G                    �?�t���?             7@=       D                    @�X�C�?
             ,@>       ?                    �?�q�q�?             @������������������������       �                     �?@       C       #             �?z�G�z�?             @A       B                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @E       F                     @      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@I       J                    �?�Q����?	             .@������������������������       �                     @K       N                     @p=
ףp�?             $@L       M       #             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @P       W                    �?     ��?
             0@Q       R                    �?x�5?,�?             "@������������������������       �                     �?S       V                    �?      �?              @T       U                    �?r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @X       Y                    �?����X�?             @������������������������       �                     @������������������������       �                      @[       ^                    �?      �?             @\       ]                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @`       g                     @x9/���?
             ,@a       f                    �?���Q��?             $@b       c       
             �?z�G�z�?             @������������������������       �                     @d       e                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @h       i       '             �?      �?             @������������������������       �                     @������������������������       �                     �?k       �                     @0`���t�?r            �g@l       �       
             �?���	�?G            �]@m       ~                    @������?            �I@n       }                    �?~�:pΈ�?             9@o       p                    �? ����?             7@������������������������       �                      @q       z                    @�&%�ݒ�?             5@r       w       !             �?.y0��k�?
             *@s       t                    �?�C��2(�?             &@������������������������       �                      @u       v                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?x       y                    �?      �?              @������������������������       �                     �?������������������������       �                     �?{       |                    �?      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                      @       �                    @���B���?             :@������������������������       �        	             3@�       �       '             �?����X�?             @������������������������       �                     @������������������������       �                      @�       �                    �?�������?)             Q@�       �       #             �?      �?              @������������������������       �                     @������������������������       �                      @�       �                    @ d��0u�?&             N@�       �                    @g_7|�?            �H@�       �                    �?����8��?            �D@�       �                    �?L36�v[�?             7@�       �                    �?      �?             0@�       �                    �?������?
             ,@�       �                    �?H�z�G�?             $@�       �                    �?      �?              @�       �                     �?؇���X�?             @������������������������       �                     @�       �       "             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                    �?؇���X�?             @������������������������       �                     @������������������������       �                     �?�       �                    @�����H�?	             2@������������������������       �                     .@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?      �?              @�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    �?��!pc�?             &@������������������������       �                     �?�       �                    @ףp=
�?             $@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    �?�� �(��?+            @Q@�       �                    �?����R�?            �D@�       �                    @�u>�?            �B@�       �                    �?R���Q�?	             4@������������������������       �                     0@�       �                    @      �?             @������������������������       �                     �?������������������������       �                     @�       �                    @�M�]��?             1@�       �                     @      �?             @������������������������       �                     �?������������������������       �                     @�       �                    @�n_Y�K�?             *@�       �                    �?      �?              @�       �       
             �?�q�q�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �       !             �?      �?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    @�r
^N��?             <@�       �                    @b�r���?             .@�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @�       �                    �?j�V���?
             &@�       �                    �?�����H�?             "@������������������������       �                     @�       �                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    �?�n_Y�K�?             *@�       �                    @z�G�z�?             $@������������������������       �                      @������������������������       �                      @������������������������       �                     @�t�bh�h)h,K ��h.��R�(KK�KK��h�B)       �A@     �E@      R@     �Y@      M@      @@      ?@      D@     �E@     �@@      @      @      &@                              @      @      $@                              @              �?                              @              �?                                                                              @              "@                                              �?                                      @      �?                                                                                      @      4@      D@     �E@     �@@                      @      .@      ,@      >@                      @       @      "@      "@                      �?      @      "@      "@                      �?      @      @                              �?       @      @                                       @      �?                                       @                                                      �?                              �?              @                              �?                                                              @                                       @                                              @      @      "@                              @      @                                       @                                              �?      @                                              @                                      �?                                                              "@                       @      �?                                       @                                                      �?                                       @      @      @      5@                       @      @                                       @      @                                              @                                       @                                                      �?                                              @      @      5@                              �?       @      5@                                              *@                              �?       @       @                              �?      �?                                              �?                                      �?                                                      �?       @                                      �?                                                       @                               @      @                                       @       @                                               @                                       @                                                      �?                              .@      9@      =@      @                      "@      5@      <@                              @      4@      <@                              @      (@      7@                               @      @      0@                               @      @      @                               @      @                                      �?                                              �?      @                                      �?      �?                                      �?                                                      �?                                              @                                              �?      @                                      �?                                                      @                                              "@                              �?      @      @                                      @                                      �?       @      @                              �?       @                                      �?                                                       @                                                      @                              @       @      @                              �?      @      @                                      �?                                      �?       @      @                              �?              @                              �?                                                              @                                       @                                       @      @                                              @                                       @                                              @      �?                                      �?      �?                                      �?                                                      �?                                       @                                              @      @      �?      @                      @      @                                      �?      @                                              @                                      �?      �?                                      �?                                                      �?                                      @                                                              �?      @                                              @                                      �?                              @      @      =@     @Q@     �K@      <@       @      @      6@      B@     �B@      3@       @      @      .@      @      5@      @       @      @      .@      @                       @      �?      .@      @                       @                                                      �?      .@      @                              �?      &@      �?                                      $@      �?                                       @                                               @      �?                                       @                                                      �?                              �?      �?                                      �?                                                      �?                                              @      @                                      @                                                      @                               @                                                                      5@      @                                      3@                                               @      @                                              @                                       @                              @      ?@      0@      ,@                               @      @                                              @                                       @                                      @      =@      $@      ,@                      @      <@      "@      @                      @      <@      @                              @      (@      @                              @      @      @                              @      @       @                              @      @      �?                              �?      @      �?                                      @      �?                                      @                                              �?      �?                                              �?                                      �?                                      �?                                               @                                              @              �?                              @                                                              �?                                               @                              �?      @                                              @                                      �?                                                      0@       @                                      .@                                              �?       @                                      �?                                                       @                                              @      @                                      @      �?                                      @                                                      �?                                              @                              �?      �?      "@                              �?                                                      �?      "@                                      �?      @                                              @                                      �?                                                      @       @              @     �@@      2@      "@                      @      9@      &@                              �?      9@      &@                                      1@      @                                      0@                                              �?      @                                      �?                                                      @                              �?       @       @                              �?      @                                      �?                                                      @                                              @       @                                      @      @                                       @      @                                      �?      �?                                              �?                                      �?                                              �?      @                                      �?      �?                                              �?                                      �?                                                       @                                       @                                              �?      @                                              @                                      �?                                      @                               @               @       @      @      "@       @               @       @       @      �?       @               @                                               @                               @                                                                       @       @      �?                               @              �?                              @                                              �?              �?                              �?                                                              �?                                       @                                              @       @                                       @       @                                       @                                                       @                                      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hKhNhJ:9)bhG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKم�h��Bx/         �                    �?�Km��?�            `u@       a                    �?���s��?�            @l@       R                    �?�j3!��?a            �d@       G                    @`.�Ň�?K            �_@       "       &             �?	|����?>            �Z@                           �?D4T2��?             G@                           �?0\�Uo��?
             3@                           �?�g���e�?             &@	                           �?������?             @
                            @      �?              @������������������������       �                     �?������������������������       �                     �?                           �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @                           @      �?              @������������������������       �                     @              #             �?      �?             @������������������������       �                     �?������������������������       �                     @                           �?<t=9%��?             ;@                           �?�"e����?             2@                           @�q�q�?             @������������������������       �                     �?������������������������       �                      @                           @�r����?             .@������������������������       �                      @������������������������       �                     *@              !             �?VUUUUU�?             "@������������������������       �                     @        !                    @      �?             @������������������������       �                     @������������������������       �                     @#       :                    @c�/��b�?%             N@$       3                    �?p@��ҽ�?             E@%       2                    �?���[���?             2@&       -                    �?     @�?             0@'       ,                     @�8��8��?             @(       +                    �?�q�q�?             @)       *                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @.       /       #             �?z�G�z�?             $@������������������������       �                     @0       1                     �?����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @4       7                    �?8��8���?             8@5       6                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?8       9                    @���N8�?             5@������������������������       �                     4@������������������������       �                     �?;       F                     �?VUUUUU�?             2@<       E                    @
ףp=
�?             $@=       >                    �?      �?              @������������������������       �                     @?       D                    �?
ףp=
�?             @@       C                    �?VUUUUU�?             @A       B                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                      @H       I                    �?�Q����?             4@������������������������       �                      @J       Q                    @VUUUUU�?	             (@K       L                    �?      �?              @������������������������       �                     @M       P       )             �?z�G�z�?             @N       O                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @S       \                    �?�P^Cy�?             C@T       W                    @J���#�?             6@U       V                    �?z�G�z�?             $@������������������������       �                      @������������������������       �                      @X       [                     @VUUUUU�?             (@Y       Z       !             �?      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     @]       ^                    @      �?
             0@������������������������       �                     &@_       `       '             �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @b       �                    �?B!�B�?.             O@c       t       %             �?,!4��=�?'            �J@d       o       !             �?x9/���?             ,@e       n       $             �?����>4�?             @f       k                    �?�8��8��?             @g       h                    �?      �?             @������������������������       �                      @i       j                    �?      �?              @������������������������       �                     �?������������������������       �                     �?l       m       "             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?p       s       '             �?0�����?             @q       r       #             �?r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?u       z                    �?x�����?            �C@v       y                    �?�$I�$I�?             @w       x                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @{       �       "             �?     ��?             @@|                           �?��ǘ���?             9@}       ~                    @8�Z$���?	             *@������������������������       �                     &@������������������������       �                      @�       �                    @9��8���?	             (@�       �                    �?      �?             @�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                    �?�q�q�?             @�       �       	             �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @�       �                    �?�$I�$I�?             @�       �                    @      �?             @������������������������       �                     �?�       �       
             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �?X�<ݚ�?             "@�       �       
             �?      �?              @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                    �?2�j�'��?E             ]@�       �                    �?�ހ2q��?5             U@�       �                    �?��e�B��?            �I@�       �                    @���}<S�?             7@������������������������       �                     2@�       �                    �?���Q��?             @������������������������       �                      @������������������������       �                     @�       �                     @@4և���?             <@������������������������       �                     1@�       �       #             �?"pc�
�?             &@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                    @�o�00s�?            �@@�       �                    �?�J�4�?             9@�       �                     �?�ӭ�a��?             2@�       �       (             �?p=
ףp�?             $@�       �       
             �?B{	�%��?             "@�       �                    �?      �?              @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    �?�$I�$I�?             @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    @      �?              @�       �                    �?�q�q�?             @������������������������       �                     �?�       �                     �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �       #             �?     @�?             @@�       �                    @��>4և�?	             ,@�       �       &             �?����X�?             @������������������������       �                      @������������������������       �                     @�       �       
             �?����X�?             @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?<ݚ)�?             2@�       �                     @޾�z�<�?             *@�       �                    �?z�G�z�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �?      �?              @������������������������       �                      @�       �                     �?�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�t�bh�h)h,K ��h.��R�(KK�KK��h�B�(        B@      P@     �U@     @R@     �O@      4@      "@      =@     @Q@      O@      H@      "@       @      8@     �M@      G@      :@      �?       @      6@     �I@      ;@      2@               @      6@     �G@      .@      ,@                      �?      5@      *@      &@                              @       @      @                              �?      @      @                              �?      @      @                              �?      �?                                      �?                                                      �?                                               @      @                                       @                                                      @                                      @                                      @      �?      @                              @                                                      �?      @                                      �?                                                      @                      �?      0@      @      @                      �?      *@       @       @                      �?               @                              �?                                                               @                                      *@               @                                               @                              *@                                              @      @      @                                      @                                      @              @                              @                                                              @               @      5@      :@       @      @              @      (@      9@      �?                      @      $@      @                              @      $@      @                              �?       @      @                              �?       @                                      �?      �?                                              �?                                      �?                                                      �?                                                      @                               @       @                                              @                                       @      @                                              @                                       @                                                               @                              �?       @      4@      �?                      �?       @                                               @                                      �?                                                              4@      �?                                      4@                                                      �?                      @      "@      �?      �?      @              @      �?      �?      �?      @               @      �?      �?      �?      @                                              @               @      �?      �?      �?                              �?      �?      �?                                      �?      �?                                      �?                                                      �?                              �?                                       @                                               @                                                       @                                                      @      (@      @                                       @                                      @      @      @                              @      @                                              @                                      @      �?                                       @      �?                                       @                                                      �?                                       @                                                              @                       @       @      3@       @      �?               @       @      @      @      �?               @       @                                       @                                                       @                                                      @      @      �?                              @              �?                                              �?                              @                                                      @                                      (@      @                                      &@                                              �?      @                                      �?                                                      @              �?      @      $@      0@      6@       @      �?      @      $@      $@      4@       @      �?      @      @      @                      �?      @      �?       @                      �?      @               @                              @              �?                               @                                              �?              �?                                              �?                              �?                                      �?                      �?                                              �?                      �?                                                              �?                                      �?      @      �?                                      @      �?                                              �?                                      @                                      �?                                                      @      @      4@       @                      @               @      �?                                       @      �?                                              �?                                       @                              @                                                      @      2@      @                              @      0@      @                                      &@       @                                      &@                                                       @                              @      @      @                              @      @                                      @      �?                                      @                                                      �?                                               @                                               @      @                                       @       @                                       @                                                       @                                               @                              @       @      �?                              �?       @      �?                              �?                                                       @      �?                                       @                                                      �?                              @                              �?              @       @                                      @       @                                      @                                              �?       @                                      �?                                                       @                      �?                                      ;@     �A@      1@      &@      .@      &@      9@      >@      0@      @      @      @      7@      <@                                      5@       @                                      2@                                              @       @                                               @                                      @                                               @      :@                                              1@                                       @      "@                                       @      �?                                              �?                                       @                                                       @                                       @       @      0@      @      @      @       @       @      0@      @                               @      .@      �?                               @      @      �?                              �?      @      �?                              �?      @                                      �?       @                                      �?                                                       @                                              @                                                      �?                              �?                                                       @                               @              �?      @                       @              �?                               @                                                              �?                                                      @                                              �?      @      @                              �?       @                                              �?                                      �?      �?                                      �?                                                      �?                                              �?      @                                              @                                      �?               @      @      �?      @      (@      @       @      @                       @      @       @      @                                       @                                                      @                                                                       @      @                                              @                                       @      �?                                       @                                                      �?                      �?      @      $@       @                      �?              $@       @                      �?              @                              �?              �?                              �?                                                              �?                                              @                                              @       @                                       @                                              @       @                                      @                                                       @                              @                �t�bubhhubh)��}�(hhhhhNhKhKhG        hKhNhJ�BHzhG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKÅ�h��B�*         �                    @1��x��?�            `u@       G       %             �?R�{�T�?�            �m@                           �?�?�0�!�?\             a@       	                    �?�g�eX�?            �A@              "             �?      �?             0@������������������������       �                     @                           @"pc�
�?             &@������������������������       �                     "@������������������������       �                      @
                           �?��N���?             3@������������������������       �                     @                            �?     ��?	             0@              
             �?���!pc�?             &@                           �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @       (                    @�g<�̉�?F            @Y@       #                    �?n�����?             B@       "                    �?�J�4�?             9@       !       $             �?������?             1@                            �?�q�q�?
             (@                           �?      �?              @                           �?      �?             @������������������������       �                      @              )             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                            �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @$       '                    �?"pc�
�?             &@%       &                    @�q�q�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                      @)       4                    �?8�w��@�?-            @P@*       /                    �?      �?             4@+       .                    �?$�q-�?             *@,       -                    �?      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     @0       1                    �?և���X�?             @������������������������       �                      @2       3                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?5       B                    �?:	��ʵ�?            �F@6       7                    �?������?            �B@������������������������       �                     0@8       9       !             �?��s����?             5@������������������������       �                     &@:       ?                    �?���Q��?             $@;       >                    �?���Q��?             @<       =                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?@       A                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @C       F                    �?      �?              @D       E                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @H       ]                    @��z��?:            @Y@I       X                    �?�S���?            �E@J       W                    �?،A��_�?
             1@K       V                    �?ƒ_,���?	             .@L       U                    �?�n_Y�K�?             *@M       P                    �?�eP*L��?             &@N       O                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?Q       R       #             �?r�q��?             @������������������������       �                      @S       T                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                      @Y       \                    �? ���c��?             :@Z       [                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     8@^       �                    @2�j�'��?#             M@_       p                    �?�q�=���?            �D@`       a       #             �?b�r���?             .@������������������������       �                      @b       m                    �?g\�5�?
             *@c       f       
             �?���(\��?             $@d       e                    �?      �?              @������������������������       �                     �?������������������������       �                     �?g       l                    �?      �?              @h       i                    �?؇���X�?             @������������������������       �                     @j       k                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?n       o                    @�q�q�?             @������������������������       �                     �?������������������������       �                      @q       v       '             �?PS!����?             :@r       u                    @      �?              @s       t                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @w       �                    �?�n����?	             2@x       }       "             �?     ��?             0@y       |                    �?8�Z$���?             *@z       {                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     "@~                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �       )             �?������?	             1@������������������������       �                     $@�       �       $             �?և���X�?             @������������������������       �                     @������������������������       �                     @�       �                    �?O��E1�??            @Z@�       �       &             �?"w|���?8            �W@�       �                    @�X�C�?)            �Q@�       �       )             �?ܤ�[r�?
             5@������������������������       �                     "@�       �                    �?�8��8��?             (@������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                    �?��eH��?            �H@�       �                    �?������?            �G@�       �                    @r��ճC�?             F@�       �                    �?�K8��?             :@�       �                    @���7�?             6@������������������������       �                     5@������������������������       �                     �?�       �                    @      �?             @������������������������       �                      @������������������������       �                      @�       �                    �?��ӭ�a�?             2@�       �                     @���Er�?             1@�       �       
             �?޾�z�<�?             *@�       �                    �?�������?             (@������������������������       �                     �?�       �                    �?�C��2(�?             &@�       �                    @z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �       	             �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    @�q�q�?             8@�       �                    �?����X�?             @������������������������       �                      @�       �                    �?���Q��?             @������������������������       �                      @�       �       !             �?�q�q�?             @������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @�IєX�?	             1@������������������������       �                     "@�       �                    �?      �?              @������������������������       �                     @������������������������       �                     �?�       �       	             �?t�E]t�?             &@�       �                    �?����>4�?             @�       �       #             �?�Q����?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @�t�bh�h)h,K ��h.��R�(KK�KK��h�B�$       �A@      J@     @V@     @R@     �P@      :@      @@      I@     @T@      B@      9@      *@      ?@      F@      G@      $@      @       @      6@       @      @                       @      ,@                                       @      @                                              "@                                       @      "@                                                                                       @       @       @      @                              @                                              @       @      @                                       @      @                                       @      @                                       @                                                      @                                      @                                      @                                              "@      B@     �E@      $@      @              @      5@      @       @      @              @      5@                                      @      *@                                      @       @                                      �?      @                                      �?      @                                               @                                      �?      �?                                      �?                                                      �?                                              @                                      @      �?                                              �?                                      @                                                      @                                               @                                                      @       @      @                              @              @                              @                                                              @                                       @                      @      .@     �B@       @                      @      .@                                      �?      (@                                      �?      @                                              @                                      �?                                                      @                                      @      @                                               @                                      @      �?                                      @                                                      �?                                                     �B@       @                                     �@@      @                                      0@                                              1@      @                                      &@                                              @      @                                       @      @                                      �?      @                                              @                                      �?                                              �?                                              @      �?                                              �?                                      @                                              @      @                                      �?      @                                      �?                                                      @                                      @                              �?      @     �A@      :@      6@      &@      �?      @      @@      @                              @       @      @                              @       @       @                              @       @                                      @      @                                      @      �?                                      @                                                      �?                                      �?      @                                               @                                      �?      @                                              @                                      �?                                                       @                                                       @                                               @                      �?      �?      8@                              �?      �?                                      �?                                                      �?                                                      8@                                              @      6@      6@      &@                      @      2@      "@      &@                       @      @      @      �?                               @                                       @      @      @      �?                      �?       @      @      �?                      �?                      �?                      �?                                                                      �?                               @      @                                      �?      @                                              @                                      �?      �?                                      �?                                                      �?                                      �?                                      �?       @                                      �?                                                       @                                      �?      (@      @      $@                      �?      �?              @                      �?      �?                                      �?                                                      �?                                                              @                              &@      @      @                              &@      @       @                              &@       @                                       @       @                                               @                                       @                                              "@                                                      �?       @                                               @                                      �?                                                       @                              @      *@                                              $@                                      @      @                                      @                                                      @              @       @       @     �B@      E@      *@      �?       @       @      >@     �D@      (@      �?              @      ,@      D@      (@                              &@      @      @                              "@                                               @      @      @                                      @                                       @              @                                              @                               @                      �?              @      @      A@       @      �?              @      @      A@      @      �?                      @      A@      @                               @      7@      �?                                      5@      �?                                      5@                                                      �?                               @       @                                       @                                                       @              �?                      �?      &@      @                              �?      &@      @                              �?      $@       @                              �?      $@      �?                              �?                                                      $@      �?                                      @      �?                                      @                                                      �?                                      @                                                      �?                                      �?      @                                      �?                                                      @      �?                                                              @                                                                       @               @      @      0@      �?                       @      @                                               @                                       @      @                                               @                                       @      �?                                      �?                                              �?      �?                                      �?                                                      �?                                                      0@      �?                                      "@                                              @      �?                                      @                                                      �?               @                      @      �?      �?       @                      @      �?      �?                              @      �?      �?                                      �?      �?                                              �?                                      �?                                      @                       @                                                                      @                �t�bub��	     hhubh)��}�(hhhhhNhKhKhG        hKhNhJ�}�JhG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK���h��B�6         �                    @4g�h�?�            `u@       s       
             �?ds�.��?�            �m@       J       )             �?�b�~wj�?[             b@       7                    �??�q�>�?7            @U@              #             �?9�b���?%             M@                           �?� ���?             ?@              !             �?�������?             4@                           �?����>4�?	             ,@	                           �?      �?              @
              %             �?      �?             @              (             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @              &             �?�q�q�?             @������������������������       �                     @                           �?�q�q�?             @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?                            @r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     &@       6       	             �?��h�C�?             ;@       )                    �?$������?             9@                            �?�8��8��?
             (@                           �?      �?             @������������������������       �                     �?������������������������       �                     @!       $                     @      �?              @"       #                     �?      �?             @������������������������       �                      @������������������������       �                      @%       (                    �?      �?             @&       '       %             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @*       5                    �?�q-�?
             *@+       4                    �?�g���e�?             &@,       3                    �?p=
ףp�?             $@-       .                    �?�<ݚ�?             "@������������������������       �                     @/       2       %             �?���Q��?             @0       1                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @8       E                    �?�ٴ��?             ;@9       @                    �?��Moz��?             7@:       ?                    �?H�z�G�?             4@;       >                    �?�d�����?             3@<       =                    �?�X�<ݺ?
             2@������������������������       �                     �?������������������������       �        	             1@������������������������       �                     �?������������������������       �                     �?A       B                     �?VUUUUU�?             @������������������������       �                     �?C       D       %             �?      �?              @������������������������       �                     �?������������������������       �                     �?F       G                    �?      �?             @������������������������       �                     �?H       I       %             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?K       R                    �?��0u���?$             N@L       M                     @:/����?             @������������������������       �                     @N       O                    �?      �?             @������������������������       �                     �?P       Q                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?S       j                    �?��M��?            �J@T       g                    �?     ��?             @@U       Z                    �?�(ݾ�z�?             :@V       Y       "             �?�<ݚ�?             "@W       X                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @[       d                    �?�hJ,��?             1@\       ]       #             �?�������?	             (@������������������������       �                     �?^       c                    @��!pc�?             &@_       `       !             �?ףp=
�?             $@������������������������       �                      @a       b                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?e       f                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @h       i                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?k       n                    �?��s����?
             5@l       m                    �?��S�ۿ?             .@������������������������       �                     ,@������������������������       �                     �?o       r       %             �?      �?             @p       q                     @���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?t       �                    �?�YY�J:�?>            �W@u       �                    �?U��6���?#            �I@v       }       %             �?����5�?             =@w       x                    �?h/�����?             "@������������������������       �                      @y       z       !             �?����X�?             @������������������������       �                      @{       |                    �?���Q��?             @������������������������       �                     @������������������������       �                      @~       �       "             �?H�z�G�?             4@       �                    �?�h$��W�?
             .@�       �                    �?�Q����?             @������������������������       �                     �?�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?�       �                    @�z�G��?             $@�       �                    �?      �?             @������������������������       �                      @�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    �?�Q����?             @������������������������       �                     �?�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �?*L�9��?             6@�       �                     �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    �?k��\��?             1@�       �                    �?�'}�'}�?             .@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �       )             �?      �?	             (@������������������������       �                     @�       �       &             �?      �?             @�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �       %             �?�ʑ���?            �E@�       �                    @      �?
             (@�       �                    �?z�G�z�?             $@������������������������       �                     @�       �                    �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @�       �                    @�����-�?             ?@�       �                    �?�ˠT��?             6@�       �                    �?�(\����?
             4@�       �                    �?�����H�?             2@�       �                    �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     *@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                     �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?�q�q�?             "@������������������������       �                     @�       �                    �?      �?             @������������������������       �                      @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?0�����?=            �Y@�       �                    @Kw�H�?$            �L@�       �       %             �?��6�K�?            �D@�       �       
             �?�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@�       �                    �?�|�j�?             >@�       �       "             �?����!p�?             6@�       �                    �?�˹�m��?             3@�       �                    @6�i�6�?             .@�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?�������?             (@�       �       )             �?�C��2(�?             &@�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?�       �                    @      �?             @������������������������       �                      @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    @     ��?
             0@�       �       %             �?r�q��?             (@������������������������       �                     �?�       �                    �?"pc�
�?             &@�       �                    �?ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?������������������������       �                     �?�       �       !             �?      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �?�ܸb���?             G@�       �                    �?����>4�?             E@�       �                    �?VUUUUU�?             .@������������������������       �                     @�       �                    �?      �?              @������������������������       �                     @�       �       !             �?      �?             @������������������������       �                     �?������������������������       �                     @�       �                    @�'��P��?             ;@�       �       !             �?�q�q�?
             5@�       �                    @�r����?             .@������������������������       �                      @������������������������       �                     *@�       �                    �?VUUUUU�?             @�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?�t�bh�h)h,K ��h.��R�(KK�KK��h�B/       �B@     @P@      N@     �U@      O@      ?@      B@     �N@     �M@      H@      6@      *@      ?@      G@     �C@      2@      @      @      :@      1@      :@      "@      @       @      7@      ,@      "@      @      @       @      1@      @      @      @               @      @      @      @      @               @      @       @      @                       @      @                                       @       @                                       @       @                                      �?       @                                                                                      �?                                              �?      @                                                       @      @                                              @                                       @      �?                                      �?      �?                                              �?                                      �?                                              �?                                              �?              @                              �?                                                              @                      &@                                              @      &@      @      �?      @              @      "@      @      �?      @              @       @      @              @              �?                              @              �?                                                                              @               @       @      @              �?               @       @                                               @                                       @                                                              @              �?                              �?              �?                              �?                                                              �?                               @                              @      @       @      �?                      @      @              �?                       @      @              �?                       @      @                                              @                                       @      @                                       @      �?                                       @                                                      �?                                               @                                                              �?                      �?                                                               @                                       @                                      @      @      1@      @      �?              �?       @      1@       @      �?                      �?      1@      �?      �?                              1@      �?      �?                              1@              �?                                              �?                              1@                                                      �?                              �?                                      �?      �?              �?                                              �?                      �?      �?                                      �?                                                      �?                                       @      �?              �?                                              �?                       @      �?                                       @                                                      �?                                      @      =@      *@      "@      �?      @      @               @                       @      @                                                               @                       @                      �?                                              �?                       @                                               @                      �?                               @      =@      &@      "@      �?      �?       @      (@      &@      @      �?      �?       @      @      $@      @      �?      �?       @      @                                       @       @                                       @                                                       @                                              @                                                      $@      @      �?      �?                      "@      �?      �?      �?                                              �?                      "@      �?      �?                              "@      �?                                       @                                              �?      �?                                              �?                                      �?                                                              �?                              �?      @                                      �?                                                      @                              @      �?                                      @                                                      �?                                      1@              @                              ,@              �?                              ,@                                                              �?                              @              @                              @               @                              @                                                               @                                              �?                      @      .@      4@      >@      0@       @      @      @      2@      &@      "@      @               @      "@       @      "@      �?               @      @       @                               @                                                      @       @                                       @                                              @       @                                      @                                                       @                                      @      @      "@      �?                      @      @       @                              �?      @      �?                                              �?                              �?      @                                              @                                      �?                                              @              @                              @              @                               @                                              �?              @                                              @                              �?                                                              @                                      @      �?      �?                                      �?                                      @              �?                              @                                                              �?      @      @      "@      @              @      �?                                      @                                              @      �?                                               @      @      "@      @                       @      �?      "@      @                       @      �?                                              �?                                       @                                                              "@      @                                      @                                              @      @                                      �?      @                                              @                                      �?                                               @                                       @                                       @      $@       @      3@      @      @       @       @               @                               @               @                              @                                              @               @                                               @                              @                                       @                                                       @       @      1@      @      @               @       @      1@      �?                       @      �?      1@                               @              0@                               @              @                                              @                               @                                                              *@                                      �?      �?                                      �?                                                      �?                                      �?              �?                                              �?                              �?                                                              @      @                                      @                                              �?      @                                               @                                      �?      �?                                      �?                                                      �?      �?      @      �?     �C@      D@      2@                      �?      =@      5@      @                      �?      :@      (@       @                              $@      �?                                              �?                                      $@                                      �?      0@      &@       @                      �?       @      &@       @                      �?      @      &@       @                      �?      @      $@      �?                      �?       @                                               @                                      �?                                                      �?      $@      �?                              �?      $@                                      �?      @                                      �?                                                      @                                              @                                                      �?                               @      �?      �?                               @                                                      �?      �?                                      �?                                                      �?                              @                                               @                                              @      "@      @                               @      "@      �?                                              �?                               @      "@                                      �?      "@                                              "@                                      �?                                              �?                                              �?              @                                              @                              �?                      �?      @              $@      3@      (@      �?      @              "@      3@      "@      �?                      @      @      @                              @                      �?                              @      @                                      @              �?                                      @      �?                                                                                      @              @               @      .@      @              @               @      .@                       @                      *@                       @                                                                      *@                       @               @       @                       @                       @                                               @                       @                                                               @                                                              @                              �?              @                                              @                              �?                �t�bubhhubh)��}�(hhhhhNhKhKhG        hKhNhJ'J�OhG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK���h��BX)         :                    �?�I�г��?�            `u@       5                    �?�Cc}h,�?@             \@                           �?Fmq��?<            �Z@                           �? �Cc}�?             <@������������������������       �        
             4@              #             �?      �?              @                            @r�q��?             @������������������������       �                     @	       
                     �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @       *                    @���5��?*            �S@       #                    �?�>4և��?             L@                           �?L紂P�?            �I@                           �?     ��?             @@              !             �?���!pc�?             6@                           �?��
ц��?             *@                           �?�q�q�?             "@                           �?���Q��?             @������������������������       �                      @������������������������       �                     @                           @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@������������������������       �                     $@              
             �?�}�+r��?             3@������������������������       �                     *@                            �?r�q��?             @������������������������       �                     @!       "                    �?      �?              @������������������������       �                     �?������������������������       �                     �?$       )                    �?���Q��?             @%       (                    �?�q�q�?             @&       '                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @+       4                    �?�X����?             6@,       -                    �?      �?
             4@������������������������       �                     @.       /                    �?�n_Y�K�?             *@������������������������       �                     @0       1                    �?      �?              @������������������������       �                     @2       3                    �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @6       9                    �?r�q��?             @7       8                    @      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @;       �                    @�5��
J�?�            �l@<       a       %             �?�-�S��?�            �h@=       F                    @��Q�^�?9             T@>       E                    @�x~fL��?            �@@?       D                    �?��!pc�?             &@@       C                    �?�q�q�?             @A       B                    �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     6@G       V                    �?���p�?#            �G@H       I                     @��a�n`�?             ?@������������������������       �                     @J       K                    �?R�}e�.�?             :@������������������������       �                     @L       O                    �?�㙢�c�?             7@M       N                    �?      �?             @������������������������       �                     @������������������������       �                     �?P       U                    @�}�+r��?             3@Q       R                    @ףp=
�?             $@������������������������       �                     @S       T                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     "@W       Z       )             �?     ��?             0@X       Y       (             �?ףp=
�?	             $@������������������������       �                     "@������������������������       �                     �?[       ^       !             �?VUUUUU�?             @\       ]                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?_       `                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?b       �                     @�g����?P            @]@c       �                    �?�q-�T�?I             Z@d       }                    �?������?9            @T@e       |                    �?dR3?т�?            �D@f       w                    �?xC�Ҁ��?            �@@g       r                    @>�Q�}�?             :@h       q                    @b�2�tk�?             2@i       p       "             �?d}h���?
             ,@j       o                    �?8�Z$���?	             *@k       l                    �?�8��8��?             (@������������������������       �                     "@m       n                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @s       t                    �?      �?              @������������������������       �                      @u       v       
             �?�q�q�?             @������������������������       �                      @������������������������       �                     @x       {                    �?0�����?             @y       z       #             �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @~       �                    �?���Q��?             D@       �                    �?�b�=y�?             9@�       �                    @9��8���?
             (@�       �                    @      �?              @�       �                     �?���Q��?             @������������������������       �                      @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �?
ц�s�?             *@�       �                    �?z�G�z�?             @�       �       )             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �       )             �?      �?              @�       �                    �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                    �?hE#߼�?
             .@�       �                    @.y0��k�?	             *@�       �                    �?�8��8��?             (@������������������������       �                      @�       �                    @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    �?������?             7@�       �                    @
ףp=
�?             .@�       �       #             �?�q�q�?             "@�       �       
             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                     @r�q��?             @������������������������       �                     �?������������������������       �                     @�       �       	             �?      �?             @������������������������       �                     @������������������������       �                     @�       �       $             �?      �?              @������������������������       �                     @������������������������       �                     �?�       �                    �?޾�z�<�?             *@������������������������       �                     $@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?����e��?            �@@�       �                    @"��u���?             9@�       �                    �?      �?             0@�       �       !             �?��S�ۿ?
             .@������������������������       �                     *@�       �                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@������������������������       �                      @�t�bh�h)h,K ��h.��R�(KK�KK��h�Bp#       �H@     �R@     �S@      R@     �I@      1@     �G@     @P@                                      E@      P@                                      9@      @                                      4@                                              @      @                                      @      �?                                      @                                               @      �?                                              �?                                       @                                                       @                                      1@     �N@                                      $@      G@                                      @      F@                                      @      :@                                      @      0@                                      @      @                                      @      @                                      @       @                                               @                                      @                                              @      �?                                      @                                                      �?                                              @                                              "@                                              $@                                      �?      2@                                              *@                                      �?      @                                              @                                      �?      �?                                              �?                                      �?                                              @       @                                      �?       @                                      �?      �?                                      �?                                                      �?                                              �?                                       @                                              @      .@                                      @      .@                                              @                                      @       @                                              @                                      @      @                                      @                                               @      @                                              @                                       @                                               @                                              @      �?                                      @      �?                                              �?                                      @                                               @                                               @      "@     �S@      R@     �I@      1@       @      "@     �S@     �Q@      =@       @       @      @     �F@      :@       @      �?       @      @      ;@                               @      @      @                               @      @                                       @      @                                       @                                                      @                                              �?                                                      @                                              6@                                              2@      :@       @      �?                      @      8@                                              @                                      @      3@                                      @                                              @      3@                                      @      �?                                      @                                                      �?                                      �?      2@                                      �?      "@                                              @                                      �?       @                                               @                                      �?                                                      "@                                      &@       @       @      �?                      "@                      �?                      "@                                                                      �?                       @       @       @                               @      �?                                       @                                                      �?                                              �?       @                                               @                                      �?                              @      A@      F@      ;@      @              @      @@      A@      :@      @              @      =@      ;@      0@      @                      3@      $@      "@      @                      &@      $@      "@      @                      &@      "@      @       @                      &@      @                                      &@      @                                      &@       @                                      &@      �?                                      "@                                               @      �?                                       @                                                      �?                                              �?                                              �?                                              @                                               @      @       @                                               @                               @      @                                       @                                                      @                                      �?      @      �?                              �?      @                                              @                                      �?                                                              �?                       @                                      @      $@      1@      @      �?              @      @      @      @      �?               @      @              @      �?               @      @               @      �?               @      @                                       @                                                      @                                                               @      �?                                      �?                                              �?      �?                                              �?                                      �?                                              @                      @      @      @                                      @      �?                                       @      �?                                              �?                                       @                                               @                                      @              @                              @               @                              @                                                               @                                              @                                      @      &@      �?                              �?      &@      �?                              �?      &@                                               @                                      �?      @                                              @                                      �?                                                              �?                               @                                              @      @      $@      @                      @      @      @      @                      @      @                                       @      �?                                       @                                                      �?                                      �?      @                                      �?                                                      @                                                      @      @                                              @                                      @                                      �?      @                                              @                                      �?                                       @      $@      �?                                      $@                                       @              �?                                              �?                               @                                                       @      6@      "@                               @      ,@      "@                               @      ,@                                      �?      ,@                                              *@                                      �?      �?                                      �?                                                      �?                                      �?                                                              "@                                       @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hKhNhJW�ehG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKͅ�h��B�,         t       
             �?l^�?�            `u@       e                    �?�3�F�?x             h@       X                    @��I.\�?f            `d@                           �?��Ku[�?]            `b@              &             �?9��8���?             8@                           �?      �?
             0@                           @؉�؉��?	             *@              !             �?ffffff�?             $@	                            @�8��8��?             @
              #             �?���Q��?             @������������������������       �                     �?                           �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @                           @      �?              @������������������������       �                     @������������������������       �                     �?       =                    �?����U+�?L            �^@       $                    �?
���?/            @R@       !       '             �?��<b���?             7@              &             �?�KM�]�?             3@������������������������       �                     �?                           �?�X�<ݺ?
             2@������������������������       �                      @                           �?ףp=
�?             $@������������������������       �                      @                             �?      �?              @������������������������       �                     �?������������������������       �                     �?"       #                     @      �?             @������������������������       �                     @������������������������       �                     �?%       &                    @�	��?!             I@������������������������       �                     $@'       8                    �?�G�z�?             D@(       7                    �?����]}�?             ;@)       6                    @�nkK�?             7@*       +                    �?�\��N��?             3@������������������������       �                      @,       -                    �?"pc�
�?             &@������������������������       �                     @.       5                    �?�q�q�?             @/       0                    �?z�G�z�?             @������������������������       �                      @1       4       %             �?�q�q�?             @2       3                     @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @9       :       #             �?8�Z$���?	             *@������������������������       �                     "@;       <       &             �?      �?             @������������������������       �                      @������������������������       �                      @>       W       	             �?/�$���?             I@?       P       %             �?�.H;T*�?            �H@@       M                    �?���?            �C@A       F       "             �?pƵHPS�?             :@B       E       !             �?և���X�?	             ,@C       D                    �?���Q��?             $@������������������������       �                     @������������������������       �                     @������������������������       �                     @G       L                    �?r�q��?             (@H       K                    @�8��8��?             @I       J                     @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @N       O                     @�	j*D�?             *@������������������������       �                     "@������������������������       �                     @Q       V                    �?���(\��?             $@R       U                    �?      �?              @S       T                    �?؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?Y       `                    @      �?	             0@Z       _                    �?      �?             $@[       \       !             �?����X�?             @������������������������       �                     �?]       ^                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @a       b                    �?r�q��?             @������������������������       �                     @c       d                    �?      �?              @������������������������       �                     �?������������������������       �                     �?f       m                    �?DDDDDD�?             >@g       l                    �?X�Cc�?
             ,@h       i       %             �?޾�z�<�?	             *@������������������������       �                     $@j       k                     �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?n       q                    �?     @�?             0@o       p                    �?r�q��?             (@������������������������       �                      @������������������������       �                     $@r       s       %             �?      �?             @������������������������       �                     @������������������������       �                     �?u       �       &             �?/�h4�p�?]            �b@v       �                    �?���M�?A             [@w       �                    @
ףp=
�?1             T@x       y       #             �?B��0�z�?            �F@������������������������       �                     .@z       �                    �?j�6�i�?             >@{       �                    �?���(\��?             4@|       �                    �?      �?
             0@}       �                    �?      �?	             (@~       �                    �?      �?              @       �                     �?      �?             @������������������������       �                      @������������������������       �                      @�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    �?p=
ףp�?             $@������������������������       �                      @�       �                    �?      �?              @������������������������       �                     @������������������������       �                     �?�       �                    �?p�_�Q�?            �A@�       �                    @�K8��?             :@�       �                    �?���7�?             6@������������������������       �                     ,@�       �                     @      �?              @������������������������       �                     @������������������������       �                     �?�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @�       �                    @h/�����?             "@�       �                    @      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    �?h�����?             <@�       �                    �?���y4F�?
             3@�       �                    �?     ��?             0@������������������������       �                      @�       �                    �?*x9/��?             ,@�       �                    @�z�G��?             $@�       �                    �?      �?             @������������������������       �                     �?�       �       #             �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �       )             �?      �?             @������������������������       �                      @������������������������       �                      @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                     @�����H�?             "@�       �                    �?z�G�z�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �?L�J��}�?            �D@�       �       $             �?�G�z��?             4@�       �       '             �?����X�?             ,@�       �                    �?      �?              @�       �                    @�q�q�?             @�       �                    �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    �?�q�q�?             5@�       �                    @�<ݚ�?             2@�       �                    @@�0�!��?             1@������������������������       �                     &@�       �                    @      �?             @�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @�t�bh�h)h,K ��h.��R�(KK�KK��h�Bp&        D@      L@     @V@     �Q@      J@      A@      =@     �E@      O@      =@      ,@      0@      0@     �C@      I@      <@      ,@      0@      0@     �C@      I@      <@       @      @      @      @       @      @      �?      @              @       @      @      �?      @              @       @      @      �?      @              @       @      @      �?                      @       @              �?                      @       @                                              �?                                      @      �?                                      @                                                      �?                                                              �?                                      @                                                              @                              @                      @                                      �?      @                                                                                      �?      "@      B@      H@      5@      @       @      @      2@      7@      5@      @              @      2@                                       @      1@                                      �?                                              �?      1@                                               @                                      �?      "@                                               @                                      �?      �?                                              �?                                      �?                                              @      �?                                      @                                                      �?                                                      7@      5@      @                              $@                                              *@      5@      @                              *@      $@      @                              "@      $@      @                              "@      $@                                               @                                      "@       @                                      @                                              @       @                                      @      �?                                       @                                               @      �?                                      �?      �?                                      �?                                                      �?                                      �?                                                      �?                                                      @                              @                                                      &@       @                                      "@                                               @       @                                       @                                                       @              @      2@      9@              �?       @      @      2@      9@              �?       @       @      2@      3@                               @      "@      .@                                       @      @                                      @      @                                      @                                                      @                                      @                                       @      �?      "@                               @      �?      @                               @      �?                                       @                                                      �?                                                      @                                              @                                      "@      @                                      "@                                                      @                              �?              @              �?       @      �?              @              �?              �?              @                                              @                              �?                                                                              �?                                                       @      �?                                                                              @      $@                                      @      @                                       @      @                                      �?                                              �?      @                                              @                                      �?                                              @                                              �?      @                                              @                                      �?      �?                                              �?                                      �?              *@      @      (@      �?                      $@      �?       @      �?                      $@               @      �?                      $@                                                               @      �?                                              �?                                       @                                      �?                                      @      @      $@                                       @      $@                                       @                                                      $@                              @      �?                                      @                                                      �?                                      &@      *@      ;@      E@      C@      2@       @       @      *@     �A@      C@      2@               @      &@     �@@      ;@      @               @      &@      >@       @                                      .@                               @      &@      .@       @                       @      $@       @                               @      @       @                               @       @       @                               @       @      @                                       @       @                                               @                                       @                                       @               @                                               @                               @                                                              @                                      @                                              @                                              �?      @       @                                               @                              �?      @                                              @                                      �?                                                      @      9@      @                              �?      7@       @                              �?      5@                                              ,@                                      �?      @                                              @                                      �?                                                       @       @                                               @                                       @                                       @       @      @                               @       @                                       @                                                       @                                                      @       @               @       @      &@      &@       @               @       @      $@      @                       @       @      "@      @                               @                                       @              "@      @                                      @      @                                      @      @                                              �?                                      @       @                                      @                                                       @                                      @                               @               @                                               @                               @                               @                              �?               @                                                                              �?                                              �?       @                                      �?      @                                      �?      �?                                              �?                                      �?                                                      @                                              @      "@      &@      ,@      @                      "@      &@                                      @      $@                                      @      @                                       @      @                                       @      @                                              @                                       @                                                      �?                                       @                                                      @                                      @      �?                                      @                                                      �?                                                      ,@      @                                      ,@      @                                      ,@      @                                      &@                                              @      @                                      �?      @                                              @                                      �?                                               @                                                      �?                                              @                �t�bub��      hhubh)��}�(hhhhhNhKhKhG        hKhNhJ���zhG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK���h��B�&         v                    @�ǂ֚:�?�            `u@       %                    �?� ���`�?�            @k@                           �?�|R���?3            �W@                           �?\�CX�?&            �Q@              "             �?z�G�z�?#            @P@                            @ףp=
�?             I@                           �?������?	             1@                           �?X�<ݚ�?             "@	       
                    @����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                      @                           �?Pa�	�?            �@@������������������������       �                     �?������������������������       �                     @@              '             �?��S���?             .@������������������������       �                     @������������������������       �                      @              
             �?      �?             @              #             �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @       $                    �?�q�q�?             8@              #             �?��S���?             .@������������������������       �                     @                           �?���|���?             &@������������������������       �                      @                            �?�<ݚ�?             "@������������������������       �                     �?        !                     @      �?              @������������������������       �                     @"       #       )             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     "@&       q                    �?��}�i9�?R            �^@'       d                     @9g�6��?H            @[@(       [                    �?��˕��?8            �S@)       F                    @����:�?/            �P@*       ?                    @<�
I��?             C@+       ,                    �?     `�?             @@������������������������       �                     �?-       <                    �?��e���?             ?@.       ;                    �?�����H�?             ;@/       4                    �?؇���X�?             5@0       1       )             �?���Q��?             @������������������������       �                      @2       3                     �?�q�q�?             @������������������������       �                      @������������������������       �                     �?5       6                    �?      �?             0@������������������������       �                     (@7       8                    �?      �?             @������������������������       �                      @9       :                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @=       >                    �?      �?             @������������������������       �                     @������������������������       �                     �?@       E                    �?      �?             @A       D                     �?      �?             @B       C                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @G       N       #             �?^N��)x�?             <@H       M                    �?�	j*D�?             *@I       J       "             �?և���X�?             @������������������������       �                      @K       L                     �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @O       Z                    �?*;L]n�?             .@P       Y                    �?�<ݚ�?             "@Q       X                    �?�$I�$I�?             @R       S                    �?      �?             @������������������������       �                     �?T       W       &             �?z�G�z�?             @U       V                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @\       a       !             �?�q�q�?	             (@]       `                    �?0�����?             @^       _                      @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @b       c                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @e       p                    @o
Z.�?             ?@f       g                    �?:���I�?
             1@������������������������       �                      @h       i                    �?hE#߼�?	             .@������������������������       �                     @j       o       !             �?x�5?,�?             "@k       n       %             �?r�q��?             @l       m                    @z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     ,@r       s                    @�X�C�?
             ,@������������������������       �                     @t       u                    �?�<ݚ�?             "@������������������������       �                      @������������������������       �                     @w       �                    @�Ȏ�W6�?P             _@x       �                    @�F�y5�?+             N@y       �                    @u�4&�o�?            �C@z       �       %             �?��)x9�?             <@{       �                    �?ܤ�[r�?             5@|       �                    �?      �?             0@}       ~                    �?~h����?             ,@������������������������       �                     @       �                    �?�g���e�?	             &@�       �                    �?�z�G��?             $@�       �                    �?      �?             @�       �       )             �?���Q��?             @�       �                    �?�q�q�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �?�$I�$I�?             @�       �                     �?      �?             @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                     @"pc�
�?	             &@������������������������       �                     @�       �                    �?      �?              @�       �                     �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                     @�E�_���?             5@������������������������       �                     �?�       �                    �?P���Q�?             4@������������������������       �                     3@������������������������       �                     �?�       �       %             �?     ��?%             P@�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @�       �                    @      �?#             N@�       �                    @���V��?            �F@������������������������       �                     C@������������������������       �                     @�       �                    �?��S���?
             .@������������������������       �                     @�       �                    �?�q�q�?             (@�       �                    @���!pc�?             &@������������������������       �                     @������������������������       �                      @������������������������       �                     �?�t�bh�h)h,K ��h.��R�(KK�KK��h�B0!        F@     @T@      K@      Q@      P@      ?@     �A@     �P@      H@      B@      2@      ,@     �@@      O@                                      0@     �K@                                      *@      J@                                      @     �F@                                      @      *@                                      @      @                                       @      @                                              @                                       @                                               @                                                       @                                      �?      @@                                      �?                                                      @@                                       @      @                                              @                                       @                                              @      @                                      �?      @                                              @                                      �?                                               @                                              1@      @                                       @      @                                      @                                              @      @                                       @                                               @      @                                      �?                                              �?      @                                              @                                      �?       @                                               @                                      �?                                              "@                                               @      @      H@      B@      2@      ,@       @      @     �E@      B@      0@      @              @      @@      3@      0@      @              @      ?@      ,@      &@      @              @      >@      @                              @      ;@      �?                              �?                                              @      ;@      �?                              @      8@                                      @      2@                                       @      @                                               @                                       @      �?                                       @                                                      �?                                      �?      .@                                              (@                                      �?      @                                               @                                      �?      �?                                      �?                                                      �?                                              @                                              @      �?                                      @                                                      �?                                      @      @                                      �?      @                                      �?      �?                                              �?                                      �?                                                       @                                       @                                              �?      $@      &@      @                                      "@      @                                      @      @                                       @                                              �?      @                                              @                                      �?                                              @                              �?      $@       @       @                      �?      @       @       @                      �?      @       @                              �?      @      �?                              �?                                                      @      �?                                      �?      �?                                      �?                                                      �?                                      @                                                      �?                                                       @                              @                                      �?      @      @      �?                              @      �?      �?                                      �?      �?                                      �?                                                      �?                              @                                      �?              @                              �?                                                              @               @      �?      &@      1@                       @      �?      &@      @                       @                                                      �?      &@      @                                      @                                      �?      @      @                              �?      @                                      �?      @                                      �?                                                      @                                              �?                                                      @                                              ,@                                      @               @      @                      @                                                               @      @                                       @                                                      @      "@      ,@      @      @@      G@      1@      "@      ,@      @      >@      �?               @      ,@      @      &@      �?               @      &@      @      @      �?              @      &@      �?      �?      �?              @      @      �?      �?      �?              @      @      �?                                      @                                      @      @      �?                              @      @                                      @      @                                      @       @                                      �?       @                                      �?      �?                                      �?                                                      �?                                              �?                                       @                                                      �?                                      @                                                              �?                                                      �?      �?                                              �?                                      �?                              @                                      �?               @      @                      �?               @      �?                                       @      �?                                       @                                                      �?                      �?                                                                      @                              @       @      @                              @                                                       @      @                                       @      �?                                              �?                                       @                                                      @                      �?              �?      3@                      �?                                                              �?      3@                                              3@                                      �?                                                       @     �F@      1@                               @               @                                               @                               @                                                     �F@      .@                                      C@      @                                      C@                                                      @                                      @       @                                      @                                              @       @                                      @       @                                      @                                                       @                                      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hKhNhJX^khG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK녔h��Bh3         p       %             �?b�����?�            `u@       I       
             �?ԦP�D�?i            �e@                           �?"�2<�t�?G            @]@                           @p=
ףp�?             $@������������������������       �                     @                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?	       @                    �?��F[~�??            �Z@
       1                    @N�jh���?7            �W@       "                    �?<'��]1�?            �H@                           �?Ua�	�?            �@@                            @P���� �?             7@                           �?�IєX�?	             1@������������������������       �                     &@                           �?r�q��?             @������������������������       �                     �?������������������������       �                     @              )             �?�q�q�?             @                           �?���Q��?             @������������������������       �                     �?              "             �?      �?             @������������������������       �                     �?                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?       !       "             �?H�z�G�?             $@                            @      �?              @������������������������       �                     @                            �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @#       $                     �?     @�?
             0@������������������������       �                     @%       .                    �?�8��8��?             (@&       -                    �?�<ݚ�?             "@'       ,                    �?������?             @(       )                    �?{�G�z�?             @������������������������       �                      @*       +       #             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                      @/       0       )             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?2       7                    �?��E���?            �F@3       4                    �?��S�ۿ?	             .@������������������������       �                     *@5       6       #             �?      �?              @������������������������       �                     �?������������������������       �                     �?8       ?       "             �?�������?             >@9       <       !             �?p�ݯ��?	             3@:       ;                    �?؇���X�?             @������������������������       �                     @������������������������       �                     �?=       >                    �?�8��8��?             (@������������������������       �                     &@������������������������       �                     �?������������������������       �                     &@A       D       !             �?*D>��?             *@B       C                    @      �?              @������������������������       �                     �?������������������������       �                     @E       F                    �?�Q����?             @������������������������       �                     @G       H                    �?      �?              @������������������������       �                     �?������������������������       �                     �?J       a                    �?������?"             L@K       ^                    �?�û��|�?             7@L       [                    �?�����?             3@M       N                    �?      �?             0@������������������������       �                     �?O       Z                    �?z�G�z�?             .@P       Y                    �?�z�G��?             $@Q       V       '             �?�<ݚ�?             "@R       S                    �?؇���X�?             @������������������������       �                     @T       U                    �?      �?              @������������������������       �                     �?������������������������       �                     �?W       X                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @\       ]                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @_       `                    �?      �?             @������������������������       �                     �?������������������������       �                     @b       o       "             �?�'�=z��?            �@@c       n                    �?��S���?             >@d       i                    �?��H�}�?             9@e       f                    @r�q��?
             2@������������������������       �                     *@g       h                    �?���Q��?             @������������������������       �                      @������������������������       �                     @j       k                    �?؇���X�?             @������������������������       �                     @l       m                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @q       �                    �?�ص�ı�?n             e@r       �       
             �?6��k�?H             [@s       �                    @pƵHP�?"             J@t       {       #             �?�f�W��?             A@u       z                    �?r�q��?             (@v       y                    �?����X�?             @w       x                     @      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     @|       �                    �?�zv�X�?             6@}       �                    �?Dy�5��?             3@~       �                    @t�E]t�?	             &@       �       '             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     @�       �                    �?      �?             @������������������������       �                     �?�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?      �?              @������������������������       �                     @�       �       '             �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    �?e������?             2@�       �                    �?؉�؉��?
             *@�       �                    @      �?              @�       �                      @�q�q�?             @������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �       !             �?z�G�z�?             @������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                    �?���Q��?             @������������������������       �                     @������������������������       �                      @�       �                    �?
^N��)�?&             L@�       �                    �?�eY�eY�?             E@�       �                    @��<�
�?            �@@�       �                    �?6�h$��?             .@�       �       #             �?�8��8��?	             (@������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?�E��ӭ�?             2@�       �                    �?�eP*L��?             &@�       �       $             �?      �?              @�       �                     �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �       (             �?h/�����?             "@�       �                    @      �?              @�       �       #             �?�q�q�?             @������������������������       �                     �?�       �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �       )             �?�m۶m��?             ,@�       �                    �?؇���X�?             @������������������������       �                     @������������������������       �                     �?�       �                    �?����X�?             @������������������������       �                     @������������������������       �                      @�       �                    @���T��?&            �N@�       �                    �?     @�?             H@�       �                    �?�n���?             "@�       �                    �?և���X�?             @������������������������       �                      @�       �       '             �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �       $             �?�^�����?            �C@�       �                    �?�eP*L��?            �@@�       �       "             �?�m۶m��?             <@�       �                    �?�G�z��?             4@�       �                    �?@4և���?	             ,@������������������������       �                     @�       �                    @      �?              @�       �       
             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    @      �?              @������������������������       �                     �?�       �                     �?և���X�?             @�       �       )             �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     @�       �                    �?8�Z$���?             *@������������������������       �                      @������������������������       �                     &@�t�bh�h)h,K ��h.��R�(KK�KK��h�B,        >@      Q@     �R@     @W@      I@      :@      9@     �N@      K@      >@       @      �?      0@     �G@      C@      *@       @      �?      @               @                      �?      @                                                               @                      �?                       @                                                                      �?      "@     �G@      B@      *@       @               @      G@      <@      $@       @              @      @@      @      @       @               @      :@      @      �?                       @      4@      �?                                      0@      �?                                      &@                                              @      �?                                              �?                                      @                                       @      @                                       @      @                                              �?                                       @       @                                      �?                                              �?       @                                      �?                                                       @                                              �?                                              @      @      �?                              @      �?      �?                              @                                                      �?      �?                                              �?                                      �?                                               @                              @      @      �?       @       @                      @                                      @       @      �?       @       @              @              �?       @       @               @              �?       @       @                              �?       @       @                                       @                                      �?               @                              �?                                                               @               @                                               @                                              �?       @                                               @                                      �?                                              �?      ,@      7@      @                      �?      ,@                                              *@                                      �?      �?                                      �?                                                      �?                                                      7@      @                                      (@      @                                      �?      @                                              @                                      �?                                              &@      �?                                      &@                                                      �?                                      &@                              �?      �?       @      @                      �?              @                              �?                                                              @                                      �?      �?      @                                              @                              �?      �?                                      �?                                                      �?                              "@      ,@      0@      1@                      "@      ,@                                      @      *@                                      @      (@                                      �?                                              @      (@                                      @      @                                       @      @                                      �?      @                                              @                                      �?      �?                                              �?                                      �?                                              �?      �?                                      �?                                                      �?                                      �?                                                      @                                       @      �?                                              �?                                       @                                              @      �?                                              �?                                      @                                                              0@      1@                                      0@      ,@                                      0@      "@                                      .@      @                                      *@                                               @      @                                       @                                                      @                                      �?      @                                              @                                      �?      �?                                              �?                                      �?                                                      @                                              @                      @      @      5@     �O@      H@      9@      @      @      2@      H@      6@       @      @      @      *@      6@      @       @      @       @      @      4@              �?                       @      $@                                       @      @                                       @       @                                       @                                                       @                                              @                                              @                      @       @      @      $@              �?      @       @      @      @              �?              �?       @      @              �?              �?       @                                               @                                      �?                                                              @              �?                              @                                              @              �?                              �?                                               @              �?                                              �?                               @                      @      �?      @                              @                                                      �?      @                                              @                                      �?                                                              @                      �?      @      @       @      @      �?      �?      �?      @       @      @      �?      �?                       @      @      �?      �?                       @                                              �?                      �?                      �?                                              �?                      �?                                                                              @      �?                                      @                                              �?      �?                                              �?                                      �?                      �?      @                                      �?                                                      @                                      @       @                                      @                                                       @                                      �?      @      :@      2@      @              �?      @      .@      0@      @              �?      �?      &@      .@      @              �?      �?      &@       @                      �?              &@                                              @                              �?              @                              �?                                                              @                                      �?               @                              �?                                                               @                                              *@      @                                      @      @                                      @       @                                       @       @                                               @                                       @                                              @                                                      @                                      @                              @      @      �?                              @      @                                      @       @                                              �?                                      @      �?                                      @                                                      �?                                               @                                                      �?                                      &@       @      �?                              @              �?                              @                                                              �?                              @       @                                      @                                                       @                              @      .@      :@      1@                      @      .@      8@      @                      @      @               @                      @      @                                       @                                              �?      @                                      �?                                                      @                                                               @                              &@      8@      @                              @      6@      @                               @      6@      @                              �?      2@      �?                              �?      *@                                              @                                      �?      @                                      �?      �?                                      �?                                                      �?                                              @                                              @      �?                                      @                                                      �?                              �?      @      @                              �?                                                      @      @                                       @      @                                       @                                                      @                                       @                                      @                                              @       @                                               @                                      @                                                       @      &@                                       @                                                      &@�t�bubhhubh)��}�(hhhhhNhKhKhG        hKhNhJQ��dhG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKӅ�h��B(.         p       
             �?��LS:�?�            `u@                           �?����3��?w             j@                           �?�F�K�P�?            �I@                           �?&L���?            �E@                           �?����K�?             B@       	       %             �?�W��H��?             A@                           @XB���?             =@������������������������       �                     <@������������������������       �                     �?
                           @�Q����?             @������������������������       �                     @                           @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                           �?�$I�$I�?             @              %             �?VUUUUU�?             @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?              "             �?      �?             @������������������������       �                     @������������������������       �                     �?                           �?      �?              @                           �?���Q��?             @������������������������       �                      @������������������������       �                     @                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?        a                    �?uT\��?Y            �c@!       4                    �?(~����?L            �`@"       -                    @F�t�K��?            �L@#       ,                    �?�r����?             >@$       +       !             �? 7���B�?             ;@%       &       '             �?�}�+r��?
             3@������������������������       �                     *@'       *                    �?r�q��?             @(       )       #             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @.       3                    �?������?             ;@/       2                    �?      �?	             ,@0       1                    �?�<ݚ�?             "@������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     *@5       T                    �?'a�����?/             S@6       M                    �?�q�1�?             H@7       J                    @{�G�z�?             D@8       G       $             �?�>���T�?            �A@9       @                    �?L]n���?             >@:       ?                    �?ףp=
�?             4@;       >                    @z�G�z�?             $@<       =       %             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     $@A       F                    �?p=
ףp�?             $@B       E                    @      �?              @C       D       (             �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                      @H       I                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @K       L                    �?���Q��?             @������������������������       �                     @������������������������       �                      @N       S                     @      �?              @O       P                    @      �?             @������������������������       �                     �?Q       R       #             �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @U       ^                    @��)x9�?             <@V       Y       %             �?���N8�?
             5@W       X                     �?      �?              @������������������������       �                     @������������������������       �                     @Z       [                    @$�q-�?             *@������������������������       �                     $@\       ]                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @_       `                    @؇���X�?             @������������������������       �                     @������������������������       �                     �?b       e                    @��8��8�?             8@c       d                    @z�G�z�?             @������������������������       �                     @������������������������       �                     �?f       o                     �?�˹�m��?
             3@g       h                    �?��Kh/�?	             2@������������������������       �                     @i       j                    �?*D>��?             *@������������������������       �                     @k       n                    �?x�5?,�?             "@l       m                     @      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?q       �                    �?˟����?Y            �`@r              %             �?�>��)��?3            @S@s       v                    �?�:m���?             >@t       u                    �?���|���?             &@������������������������       �                     @������������������������       �                     @w       ~                    @p�ݯ��?             3@x       {                    �?؇���X�?	             ,@y       z                    �?�8��8��?             (@������������������������       �                     &@������������������������       �                     �?|       }                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    @�%��-�?             �G@�       �       $             �?�L:�d�?            �@@�       �                    �?9��8���?             8@�       �                    @ףp=
��?             4@�       �                    @      �?              @�       �                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?�       �       )             �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?�q�q�?
             (@������������������������       �                     �?�       �                    �?���!pc�?	             &@�       �       #             �?r�q��?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    @���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                    @B{	�%��?             "@�       �                     @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �       "             �?T�r
^N�?             ,@�       �                    �?���!pc�?             &@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?V��_���?&            �L@�       �                    @d���q�?            �D@�       �       %             �?b���i��?             &@�       �                    �?z�G�z�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                     �?      �?             @������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @hE#߼�?             >@������������������������       �                     @�       �                    @.y0��k�?             :@�       �                    �?�C��2(�?             6@�       �                    �?P���Q�?             4@������������������������       �                     (@�       �                    @      �?              @�       �                     @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    @      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @      �?             @������������������������       �                      @������������������������       �                      @�       �                    �?     @�?             0@�       �                    �?�g���e�?             &@�       �       %             �?�z�G��?             $@������������������������       �                     �?�       �                    �?�<ݚ�?             "@������������������������       �                     �?�       �                    @      �?              @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                    @{�G�z�?             @������������������������       �                     �?�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @�t�bh�h)h,K ��h.��R�(KK�KK��h�B�'        H@     �P@     �Q@      S@      J@      <@     �D@      L@      G@      ?@      7@      &@      >@      @      $@      @      @       @      >@      �?      @      �?      @      �?      <@              @      �?      @      �?      <@              @      �?      �?      �?      <@                      �?                      <@                                                                      �?                                      @              �?      �?                      @                                                              �?      �?                                      �?                                                      �?                                       @               @      �?      @                              �?      �?      �?                              �?              �?                              �?                                                              �?                                      �?                                      �?              @                                              @                              �?                                                       @      @       @              �?               @      @                                       @                                                      @                                                       @              �?                               @                                                              �?      &@     �J@      B@      <@      4@      "@      &@      J@      ?@      ;@      $@       @      &@      G@                                      @      :@                                      �?      :@                                      �?      2@                                              *@                                      �?      @                                      �?      �?                                      �?                                                      �?                                              @                                               @                                      @                                              @      4@                                      @      @                                       @      @                                              @                                       @                                              @                                                      *@                                              @      ?@      ;@      $@       @              @      :@      &@      @      �?              @      :@       @                              @      :@      @                              @      9@       @                               @      2@                                       @       @                                       @      �?                                       @                                                      �?                                              @                                              $@                                      �?      @       @                              �?      @                                      �?      @                                              @                                      �?                                                      @                                                       @                                      �?      @                                      �?                                                      @                              @               @                              @                                                               @                                              @      @      �?                              �?      @      �?                              �?                                                      @      �?                                              �?                                      @                                       @                                      @      0@      @      �?                      @      0@                                      @      @                                              @                                      @                                              �?      (@                                              $@                                      �?       @                                      �?                                                       @                                                      @      �?                                      @                                                      �?              �?      @      �?      $@      @                      @      �?                                      @                                                      �?                              �?      �?              $@      @                      �?              $@      @                                      @                              �?              @      @                                              @                      �?              @      @                                      @      @                                      @                                                      @                      �?                                      �?                                      @      &@      9@     �F@      =@      1@      @      @      3@      3@      7@      @      @      @      (@      @                      @      @                                              @                                      @                                                              (@      @                                      (@       @                                      &@      �?                                      &@                                                      �?                                      �?      �?                                              �?                                      �?                                                      @                                      @      (@      7@      @                      @      &@      .@                              @      $@       @                              @      $@      @                              @       @                                      @      �?                                      @                                                      �?                                      �?      �?                                      �?                                                      �?                                               @      @                                              �?                                       @      @                                      @      �?                                      �?      �?                                              �?                                      �?                                              @                                              @       @                                      @                                                       @                                              @                              �?      �?      @                              �?      �?                                      �?                                                      �?                                                      @                                      �?       @      @                                       @      @                                      �?      @                                              @                                      �?                                              @                                      �?               @                                               @                              �?                      @      @      @      :@      @      (@      �?      @      @      7@      @      @      �?      @              �?      �?      @      �?      @                                      �?      �?                                      �?                                                      �?                                              @                                                              �?      �?      @                                              @                              �?      �?                                      �?                                                      �?                              @      6@       @                              @                                               @      6@       @                               @      4@                                      �?      3@                                              (@                                      �?      @                                      �?       @                                      �?                                                       @                                              @                                      �?      �?                                              �?                                      �?                                                       @       @                                       @                                                       @               @                      @      @       @                              @      �?      @                              @              @                              �?                                               @              @                              �?                                              �?              @                              �?               @                              �?                                                               @                                              @                                      �?               @                               @      �?                                              �?       @                               @               @                                                                               @        �t�bub��     hhubh)��}�(hhhhhNhKhKhG        hKhNhJ���lhG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK���h��Bh%         P       %             �?���,Q�?�            `u@       '                    �?���`5�?j            @d@                           �?,ZYN(��?8            @T@                            �?�KM�]�?
             3@                           �?����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     (@	                           �?j�g�y�?.             O@
                           �?*
;&���?!             G@              	             �?�}�+r��?             3@������������������������       �                     1@                           �?      �?              @������������������������       �                     �?������������������������       �                     �?                           �?�<ݚ�?             ;@                           �?$�q-�?             *@������������������������       �                     (@������������������������       �                     �?                           �?X�Cc�?             ,@                           @      �?             @������������������������       �                     @������������������������       �                     �?                           �?z�G�z�?             $@              "             �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @                            �?      �?             0@                            �?؇���X�?             @������������������������       �                     �?������������������������       �                     @!       "                      @�<ݚ�?             "@������������������������       �                     @#       &       )             �?�q�q�?             @$       %                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @(       A                    �?��޸���?2            @T@)       0                    �?e������?             B@*       /                    �?      �?              @+       .       (             �?z�G�z�?             @,       -                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @1       6                    @���>4��?             <@2       3                     @VUUUUU�?             @������������������������       �                      @4       5                    �?      �?             @������������������������       �                      @������������������������       �                      @7       <                    �?��2(&�?             6@8       9                    @      �?             0@������������������������       �                     (@:       ;                     �?      �?             @������������������������       �                     @������������������������       �                     �?=       >       '             �?�q�q�?             @������������������������       �                     @?       @       
             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?B       E                    @��㜏�?            �F@C       D                    �?@4և���?             ,@������������������������       �                     �?������������������������       �                     *@F       O                    �?��a�n`�?             ?@G       N       
             �?�X����?             6@H       M                    �?���|���?             &@I       J       #             �?      �?              @������������������������       �                     @K       L                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     &@������������������������       �                     "@Q       �                    @���=�?q            �f@R       ]                    @e��z�?;            �W@S       X                    �?6�����?             5@T       W                    �?     ��?	             0@U       V       #             �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     (@Y       \       '             �?�Q����?             @Z       [                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @^       e                    �?�i��^�?/            @R@_       d                     �?��Q��?             $@`       c                    @{�G�z�?             @a       b                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @f                           �?L�!�V��?)            �O@g       ~                    �?�o�u<��?            �D@h       {                    �?pB躍�?             A@i       n                    �?�o_��?             9@j       m       !             �?      �?              @k       l                      @���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @o       z                     @��\���?             1@p       u       
             �?�������?             (@q       t                    �?�q�q�?             @r       s                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?v       y       '             �?�����H�?             "@w       x                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @|       }                    �?�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �?���7�?             6@������������������������       �                     3@�       �                    �?�q�q�?             @������������������������       �                     �?�       �                    @      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @�QK���?6            �U@�       �                    �?�{��?��?"             K@�       �                    �?J�8���?             =@�       �                    @      �?             8@�       �       !             �?և���X�?	             ,@�       �                    �?���!pc�?             &@�       �                    �?z�G�z�?             $@�       �       (             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �        	             $@�       �                    @z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    �?`2U0*��?             9@������������������������       �                     8@������������������������       �                     �?�       �       	             �?      �?             @@�       �                    �?�LQ�1	�?             7@�       �       )             �?��S���?             .@�       �                    �?      �?              @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     �?�       �       (             �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @؇���X�?             @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     "@�t�bh�h)h,K ��h.��R�(KK�KK��h�B        �D@     �L@     @R@      V@     �K@      <@     �A@      J@      D@      =@       @      @      @@     �H@                                      1@       @                                      @       @                                      @                                                       @                                      (@                                              .@     �G@                                      @     �C@                                      �?      2@                                              1@                                      �?      �?                                      �?                                                      �?                                      @      5@                                      �?      (@                                              (@                                      �?                                              @      "@                                      @      �?                                      @                                                      �?                                       @       @                                       @      @                                              @                                       @                                                      @                                       @       @                                      @      �?                                              �?                                      @                                               @      @                                              @                                       @      @                                       @      �?                                       @                                                      �?                                              @                                      @      @      D@      =@       @      @      @       @      4@      @       @      @      @              �?                      @                      �?                      @                      �?                       @                                               @                      �?                                                                       @      @                                                       @      3@      @       @                       @               @       @                       @                                                               @       @                                               @                                       @                                      3@      @                                      .@      �?                                      (@                                              @      �?                                      @                                                      �?                                      @       @                                      @                                              �?       @                                               @                                      �?                                      �?      4@      8@                              �?      *@                                      �?                                                      *@                                              @      8@                                      @      .@                                      @      @                                      @      �?                                      @                                              @      �?                                      @                                                      �?                                              @                                              &@                                              "@                      @      @     �@@     �M@     �J@      8@      @      @     �@@      H@       @              @       @      *@                              @      �?      (@                              @      �?                                      @                                                      �?                                                      (@                              @      �?      �?                                      �?      �?                                              �?                                      �?                                      @                                                      @      4@      H@       @                       @      @      �?       @                       @              �?       @                       @              �?                                              �?                               @                                                                       @                              @                                      �?      .@     �G@                              �?      ,@      :@                              �?      ,@      3@                              �?      *@      &@                                      @      @                                      @       @                                               @                                      @                                                      @                              �?      $@      @                              �?      $@      �?                              �?       @                                      �?      �?                                      �?                                                      �?                                              �?                                               @      �?                                       @      �?                                       @                                                      �?                                      @                                                      @                                      �?       @                                               @                                      �?                                                      @                                      �?      5@                                              3@                                      �?       @                                              �?                                      �?      �?                                              �?                                      �?                                                      &@     �I@      8@                              &@     �E@                                      $@      3@                                      @      2@                                      @       @                                      @       @                                       @       @                                       @      �?                                              �?                                       @                                                      @                                      �?                                              @                                                      $@                                      @      �?                                      @                                                      �?                                      �?      8@                                              8@                                      �?                                                       @      8@                                       @      .@                                       @      @                                      @      �?                                      @                                               @      �?                                      �?                                              �?      �?                                              �?                                      �?                                              �?      @                                              @                                      �?       @                                      �?                                                       @                                               @                                              "@�t�bubhhubh)��}�(hhhhhNhKhKhG        hKhNhJB	VhG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKǅ�h��B�+         b       %             �?��c����?�            `u@       W                    �?͎Z���?o             e@                           �?x�Q���?h             c@              (             �?^s]ev�?             =@                           �?�6|����?             :@              #             �?�J�4�?             9@       
                     �?      �?             0@       	                    �?      �?             @������������������������       �                      @������������������������       �                      @                           �?r�q��?
             (@              $             �?      �?              @������������������������       �                     @                           @      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     "@������������������������       �                     �?������������������������       �                     @       ,                    �?�rT���?S             _@       +                    �?F�4�Dj�?#            �M@       *       	             �?��|�5��?            �G@       )                     �?�T|n�q�?            �E@       $                    @     ��?             @@       #       "             �?R���Q�?             4@                           �?�KM�]�?             3@������������������������       �                     $@       "                    �?�<ݚ�?             "@       !                    �?      �?              @                            �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     �?%       (       !             �?�q�q�?             (@&       '                    �?և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     &@������������������������       �                     @������������������������       �                     (@-       2                    �?`�S^o�?0            @P@.       1       (             �?{�G�z�?             @/       0                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @3       N       
             �?�gE#��?-             N@4       M       "             �?*�8�G��?             A@5       L       (             �?���QI�?             9@6       K                    @�������?             8@7       H                    @���x�?             7@8       9       !             �?p=
ףp�?             4@������������������������       �                      @:       ?                    �?�q�q�?
             (@;       <                    �?r�q��?             @������������������������       �                     @=       >       )             �?      �?              @������������������������       �                     �?������������������������       �                     �?@       G                    �?      �?             @A       F       $             �?���Q��?             @B       E                    �?      �?             @C       D                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     �?I       J                    @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@O       V                    @$��m��?             :@P       U                    �?      �?             (@Q       T                    �?"pc�
�?
             &@R       S                    @ףp=
�?	             $@������������������������       �                     "@������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �        	             ,@X       _                    �?��A���?             .@Y       Z                    �?r�q��?             (@������������������������       �                      @[       ^                     @ףp=
�?             $@\       ]                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @`       a                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?c       �                    @��ys�?q            �e@d       m                    �?B�0�~��?:             V@e       j       
             �?     ��?	             0@f       g                    �?؇���X�?             ,@������������������������       �                      @h       i                    �?�q�q�?             @������������������������       �                      @������������������������       �                     @k       l                    �?      �?              @������������������������       �                     �?������������������������       �                     �?n       �       !             �?�Hx�5�?1             R@o       �                    @J���#��?!             F@p       q                    @�o_��?             9@������������������������       �                     @r              "             �?<ݚ)�?             2@s       t                    @��A���?             .@������������������������       �                     @u       v                    @{�G�z�?             $@������������������������       �                     �?w       ~                     �?x�5?,�?             "@x       {       
             �?�8��8��?             @y       z                    �?      �?              @������������������������       �                     �?������������������������       �                     �?|       }                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �?�lO���?             3@�       �       
             �?�����H�?             2@�       �                    �?z�G�z�?             $@������������������������       �                     �?�       �                    @�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                    �?ܶm۶m�?             <@������������������������       �                     (@�       �                    �?     ��?
             0@������������������������       �                      @�       �                    �?�m۶m��?             ,@�       �                    �?8�Z$���?             *@������������������������       �                     &@������������������������       �                      @������������������������       �                     �?�       �                    �?r�lUO��?7            �U@�       �                    �?����7�?/            @S@�       �                    �?؇���X�?             @������������������������       �                     @�       �       "             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?p�_�Q�?+            �Q@�       �                    @�lO���?             C@�       �                    �?(N:!���?            �A@�       �       "             �?�FVQ&�?            �@@�       �                     @�g�y��?             ?@������������������������       �                     <@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �       !             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                     �?     @�?             @@�       �                    @�����H�?             "@������������������������       �                      @������������������������       �                     �?�       �                    @�㙢�c�?             7@�       �                    �?�$I�$I�?
             ,@�       �                    @      �?	             (@������������������������       �                      @�       �       )             �?z�G�z�?             $@������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �       	             �?�<ݚ�?             "@�       �       '             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �       $             �?�n���?             "@�       �                    �?{�G�z�?             @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?�t�bh�h)h,K ��h.��R�(KK�KK��h�BP%        A@      M@     �T@     @T@     �M@      ;@     �@@      K@      I@      7@      @      @      @@     �J@     �D@      5@      @      @      5@      @      @      �?                      5@              @      �?                      5@              @                              (@              @                               @               @                               @                                                               @                              $@               @                              @               @                              @                                               @               @                               @                                                               @                              @                                              "@                                                                      �?                              @                                      &@      I@     �B@      4@      @      @      &@      H@                                      &@      B@                                      @      B@                                      @      9@                                      @      1@                                       @      1@                                              $@                                       @      @                                      �?      @                                      �?      @                                              @                                      �?                                                      @                                      �?                                              �?                                              @       @                                      @      @                                      @                                                      @                                              @                                              &@                                      @                                                      (@                                               @     �B@      4@      @      @                      �?               @       @                      �?               @                                               @                              �?                                                                       @               @      B@      4@      �?      �?               @      ;@      @      �?      �?               @      2@      @      �?      �?              �?      2@      @      �?      �?              �?      2@      @      �?                      �?      0@      @                                       @                                      �?       @      @                              �?      @                                              @                                      �?      �?                                              �?                                      �?                                                      @      @                                       @      @                                      �?      @                                      �?      �?                                              �?                                      �?                                                       @                                      �?                                              �?                                               @              �?                                              �?                               @                                                                      �?              �?                                                      "@                                              "@      1@                                      "@      @                                      "@       @                                      "@      �?                                      "@                                                      �?                                              �?                                              �?                                              ,@                      �?      �?      "@       @               @              �?      "@                       @                                               @              �?      "@                                      �?       @                                      �?                                                       @                                              @                              �?                       @                                               @                      �?                                              �?      @     �@@      M@      L@      6@      �?      @     �@@      H@       @                       @      (@      �?      �?                       @      (@                                               @                                       @      @                                       @                                                      @                                                      �?      �?                                              �?                                      �?                      �?       @      5@     �G@      �?              �?      �?      1@      8@      �?              �?      �?      .@       @                                      @                              �?      �?       @       @                      �?      �?       @      @                                      @                              �?      �?      @      @                              �?                                      �?              @      @                      �?              @       @                      �?                      �?                                              �?                      �?                                                              @      �?                                      @                                                      �?                                              @                                              @                                       @      0@      �?                               @      0@                                       @       @                                      �?                                              �?       @                                               @                                      �?                                                       @                                                      �?                      �?      @      7@                                              (@                              �?      @      &@                                       @                                      �?       @      &@                                       @      &@                                              &@                                       @                                      �?                                                              $@      K@      6@                              @     �I@      4@                                      �?      @                                              @                                      �?       @                                               @                                      �?                                      @      I@      ,@                              @      @@       @                              @      ?@                                       @      ?@                                      �?      >@                                              <@                                      �?       @                                      �?                                                       @                                      �?      �?                                      �?                                                      �?                                       @                                                      �?       @                                               @                                      �?                                       @      2@      (@                                       @      �?                                       @                                                      �?                               @      $@      &@                               @       @      @                               @       @       @                               @                                                       @       @                                      @                                              �?       @                                      �?                                                       @                                               @                                       @      @                                       @      �?                                              �?                                       @                                                      @                              @      @       @                              �?       @       @                                      �?       @                                               @                                      �?                                      �?      �?                                      �?                                                      �?                                      @      �?                                      @                                                      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hKhNhJMk/hG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKх�h��B�-         j       &             �?�*���?�            `u@       E                    @,2��.�?t            �f@       D       "             �?vSAٴ�?=            @W@       /                    �?���$�?5            �T@       .                    @I�$I�$�?#             L@       -                    �?�������?             H@                           �?ɶ���?            �C@                           �?      �?              @	       
                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @                           �?��rT��?             ?@                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?       ,                     @�m۶m��?             <@              #             �?Έ����?             9@                           �?�$I�$I�?             @������������������������       �                     @                           �?      �?             @������������������������       �                      @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?       +                    �?�[��"e�?             2@               
             �?     ��?             0@                           �?r�q��?             @������������������������       �                     @                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @!       *                    �?���Q��?             $@"       #                    �?�q�q�?             "@������������������������       �                     @$       )       '             �?      �?             @%       &                    �?���Q��?             @������������������������       �                      @'       (                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     "@������������������������       �                      @0       3       #             �?��WV��?             :@1       2                    �?�q�q�?             @������������������������       �                      @������������������������       �                     @4       ;                    �?p=
ףp�?             4@5       6                     @:/����?             @������������������������       �                      @7       :                     �?���Q��?             @8       9                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @<       C                    @8�Z$���?	             *@=       >                    �?���Q��?             @������������������������       �                      @?       @       '             �?�q�q�?             @������������������������       �                     �?A       B                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     &@F       c                    �?�L��7Q�?7            @V@G       `                    @<�;��?/            �S@H       Y                    @�p�F�:�?(            @Q@I       X                    �?�g���e�?             6@J       W       (             �?և���X�?             5@K       P                    �?(������?             3@L       O                    �?r�q��?             (@M       N                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     "@Q       R       #             �?և���X�?             @������������������������       �                     �?S       T                     @      �?             @������������������������       �                      @U       V                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?Z       [                    �?��0{9�?            �G@������������������������       �                     9@\       ]                    @�X����?             6@������������������������       �                     @^       _                    @     ��?
             0@������������������������       �                     "@������������������������       �                     @a       b                    @�q�q�?             "@������������������������       �                     @������������������������       �                     @d       i                     �?��ˠ�?             &@e       h                    �?������?             @f       g                    @      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     @k       �                    �?��(\���?f             d@l       �       #             �?.F.@�;�?U             `@m       �                    �? �2,?��?&            �M@n       �                    �?�琚`��?"            �J@o       r                    �?l �&��?             G@p       q                    �?      �?             @������������������������       �                     @������������������������       �                     @s       �       !             �?�z�G��?             D@t       {                    @g\�5�?             :@u       x                    �?�$I�$I�?             @v       w                     @�q�q�?             @������������������������       �                      @������������������������       �                     �?y       z                    �?      �?             @������������������������       �                     @������������������������       �                     �?|       �                    �?�d�����?	             3@}       �                      @�IєX�?             1@~                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     ,@�       �       "             �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?���>4��?
             ,@�       �                     @������?             @������������������������       �                     @�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �?������?             @�       �       "             �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    �?������?             @�       �                     @      �?             @������������������������       �                     �?������������������������       �                     @�       �                    @�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                     @r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                    �?����:�?/            �Q@�       �                    �?tk~X��?             B@�       �                    �?     ��?             @@�       �       !             �?      �?             8@�       �                    �?     ��?
             0@�       �                     �?@4և���?             ,@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@������������������������       �                      @������������������������       �                      @�       �                    �?      �?              @�       �                    �?�q�q�?             @�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    @�E��'s�?             A@�       �                    �?���Y �?             ;@�       �                    @�6|����?             :@�       �                    �?���}<S�?             7@������������������������       �                     *@�       �                    @z�G�z�?	             $@������������������������       �                     @�       �                    �?���Q��?             @������������������������       �                     @������������������������       �                      @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                    �?؇���X�?             @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �       !             �?�����?             ?@�       �                    �?��u0f��?             ;@�       �                     @>W[����?             9@�       �                    �?�GN�z�?             6@�       �                    @      �?	             0@������������������������       �                     $@�       �                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �       )             �?      �?             @������������������������       �                     @������������������������       �                     �?�t�bh�h)h,K ��h.��R�(KK�KK��h�B0'       �B@      H@      W@     �S@     @P@      5@      �?      @      C@     �L@      P@      2@      �?      @      C@      G@      @              �?      @      C@     �A@      @              �?      @      >@      5@                      �?      @      >@      *@                      �?      @      5@      *@                              �?      @                                      �?      @                                              @                                      �?                                                      @                              �?      @      ,@      *@                      �?               @                                               @                              �?                                                      @      (@      *@                              @      (@      $@                               @      �?      @                                              @                               @      �?      �?                               @                                                      �?      �?                                              �?                                      �?                                      �?      &@      @                              �?      &@      @                              �?      @                                              @                                      �?       @                                      �?                                                       @                                              @      @                                      @      @                                      @                                              @      @                                       @      @                                               @                                       @      �?                                       @                                                      �?                                      �?                                                      �?                                               @                                              @                                      "@                                                       @                                       @      ,@      @                              @               @                                               @                              @                                              @      ,@       @                               @      @       @                                               @                               @      @                                       @      �?                                       @                                                      �?                                               @                                       @      &@                                       @      @                                               @                                       @      �?                                      �?                                              �?      �?                                              �?                                      �?                                                       @                                              &@                                              &@      N@      2@                              @     �L@      .@                              @      K@      "@                              @      ,@       @                              @      ,@       @                              @      ,@       @                                      $@       @                                      �?       @                                      �?                                                       @                                      "@                                      @      @                                              �?                                      @      @                                               @                                      @      �?                                      @                                                      �?                                       @                                              �?                                                      D@      @                                      9@                                              .@      @                                      @                                              "@      @                                      "@                                                      @                                      @      @                                      @                                                      @                              @      @      @                              �?      @      @                                      @      @                                              @                                      @                                      �?                                              @                      B@      F@      K@      6@      �?      @      2@     �C@      H@      4@      �?      @      &@      $@      :@      "@              @      $@      $@      :@      @              @      @      @      9@      @              @      @                                      @                                              @      @                                              @      @      9@      @                      �?      @      5@      �?                      �?       @      @                                       @      �?                                       @                                                      �?                              �?              @                                              @                              �?                                                      �?      1@      �?                              �?      0@                                      �?       @                                               @                                      �?                                                      ,@                                              �?      �?                                      �?                                                      �?                      @      @      @      @                              @      �?      @                              @                                                      �?      @                                      �?                                                      @                      @      �?      @                              @      �?                                      @                                                      �?                                                      @                              @      @      �?                              �?      @                                      �?                                                      @                                       @              �?                                              �?                               @                                              �?                      @                      �?                                                                      @                      @      =@      6@      &@      �?              @      =@                                      @      9@                                      @      5@                                      @      *@                                      �?      *@                                      �?      �?                                      �?                                                      �?                                              (@                                       @                                                       @                                      @      @                                      @       @                                      @      �?                                              �?                                      @                                                      �?                                               @                                              @                                                      6@      &@      �?                              5@      @      �?                              5@      @      �?                              5@       @                                      *@                                               @       @                                      @                                              @       @                                      @                                                       @                                               @      �?                                              �?                                       @                                              �?                                      �?      @                                              @                                      �?       @                                      �?                                                       @                      2@      @      @       @                      1@      @      @       @                      1@      @      @                              1@      @                                      .@      �?                                      $@                                              @      �?                                      @                                                      �?                                       @      @                                       @                                                      @                                                      @                                                       @                      �?              @                                              @                              �?                                        �t�bubhhubh)��}�(hhhhhNhKhKhG        hKhNhJH�_VhG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK���h��B�'         .                    �?^$����?�            `u@                           �?���o_�?;             Y@                           �?6YE�t�?            �@@������������������������       �                     5@                           �?�q�q�?             (@              !             �?      �?              @              &             �?����X�?             @������������������������       �                      @	       
                    �?���Q��?             @������������������������       �                      @              )             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @                           �?��ga�=�?'            �P@                            @ܷ��?��?             =@������������������������       �                     &@                            �?r�q��?
             2@                           �?@4և���?             ,@������������������������       �                     �?������������������������       �                     *@              "             �?      �?             @                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?       -                    �?�����?             C@       *       
             �?և���X�?             <@       )                    �?������?             1@       $                    �?���|���?             &@        #                    �?؇���X�?             @!       "                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @%       (                    �?      �?             @&       '                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @+       ,                    �?���!pc�?             &@������������������������       �                     @������������������������       �                      @������������������������       �                     $@/       �                    @�H�}���?�            @n@0       y                    @�B�B1�?T            �^@1       x                    @�a�H�/�?F            �Y@2       Y                    �?�s����?E             Y@3       F                    @�i�qK�?/            �Q@4       ?                    �?      �?              H@5       <                    �?����[��?             B@6       ;                    @(;L]n�?             >@7       8                     @�8��8��?	             (@������������������������       �                     $@9       :                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     2@=       >                    �?�q�q�?             @������������������������       �                     @������������������������       �                      @@       C                    �?r�q��?	             (@A       B                     �?�����H�?             "@������������������������       �                      @������������������������       �                     �?D       E       )             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @G       T                     @�zv�X�?             6@H       Q                    �?��>4և�?	             ,@I       N                    �?��E���?             "@J       M                    �?r�q��?             @K       L       #             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @O       P       
             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?R       S                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?U       X                    �?      �?              @V       W       
             �?r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @Z       m                    �?�q�q�?             >@[       j                    �? )O��?             2@\       g       (             �?     @�?             0@]       d       
             �?*D>��?
             *@^       c                    �?B{	�%��?             "@_       b                    �?      �?              @`       a                     �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?e       f                    �?      �?             @������������������������       �                     @������������������������       �                     �?h       i                    @�q�q�?             @������������������������       �                     �?������������������������       �                      @k       l                    �?      �?              @������������������������       �                     �?������������������������       �                     �?n       w                    �?��8��8�?             (@o       p                    �?�z�G��?             $@������������������������       �                     @q       v                    �?���Q��?             @r       s       '             �?      �?             @������������������������       �                      @t       u                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @z       {                    @�Q����?             4@������������������������       �                     @|       }                    �?�t����?             1@������������������������       �                     *@~                           �?      �?             @������������������������       �                      @������������������������       �                      @�       �                    @:m���?G             ^@�       �                    �?]��$E�?0            @T@�       �                     @���
l�?)            �Q@�       �                    @     ��?'             P@�       �       
             �?>��C��?            �E@�       �                    @�z�G��?	             $@�       �                    �?      �?             @�       �                    �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    �?�C��2(�?            �@@�       �                    �?      �?             (@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     5@�       �                    �?�����?             5@������������������������       �                     3@������������������������       �                      @�       �                    @�q�q�?             @������������������������       �                     @������������������������       �                      @�       �       %             �?j�V���?             &@������������������������       �                     @�       �                    �?      �?             @������������������������       �                      @�       �       )             �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?j]%B���?            �C@�       �                    �?t���?             7@�       �       
             �?�IєX�?             1@�       �       '             �?z�G�z�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     (@�       �                    �?�8��8��?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @      �?             @������������������������       �                     @������������������������       �                     �?�       �                    @     ��?	             0@������������������������       �                     @�       �                    @�z�G��?             $@������������������������       �                     @������������������������       �                     @�t�b�8     h�h)h,K ��h.��R�(KK�KK��h�B�!        F@      N@      U@     �S@     �N@      .@     �E@     �L@                                      <@      @                                      5@                                              @      @                                      @      @                                       @      @                                               @                                       @      @                                               @                                       @      �?                                              �?                                       @                                              �?                                              @                                              .@      J@                                      @      :@                                              &@                                      @      .@                                      �?      *@                                      �?                                                      *@                                       @       @                                      �?       @                                               @                                      �?                                              �?                                              (@      :@                                      (@      0@                                      @      *@                                      @      @                                      �?      @                                      �?      @                                              @                                      �?                                                      @                                      @      �?                                       @      �?                                              �?                                       @                                              �?                                                      @                                       @      @                                              @                                       @                                                      $@                                      �?      @      U@     �S@     �N@      .@      �?      @      O@      C@      *@      @      �?      @     �M@      7@      &@      @      �?      @     �M@      7@      "@      @      �?      �?      H@      *@      @       @      �?      �?      E@      @                              �?     �@@       @                              �?      =@                                      �?      &@                                              $@                                      �?      �?                                      �?                                                      �?                                              2@                                              @       @                                      @                                                       @                      �?              "@       @                      �?               @                                               @                              �?                                                              �?       @                                      �?                                                       @                                      @      "@      @       @                      @       @      @       @                      �?      �?      @       @                      �?              @                              �?              �?                                              �?                              �?                                                              @                                      �?               @                                               @                              �?                                      @      �?                                      @                                                      �?                                      �?      @                                      �?      @                                      �?                                                      @                                               @                               @      &@      $@      @      @               @       @      @      @      �?               @       @      @      @                      �?       @      �?      @                      �?      @      �?                              �?      @                                      �?       @                                      �?                                                       @                                              @                                                      �?                                      �?              @                                              @                              �?                                      �?               @                              �?                                                               @                                                      �?      �?                                              �?                                      �?                              @      @               @                      @      @                                              @                                      @       @                                      @      �?                                       @                                              �?      �?                                      �?                                                      �?                                              �?                                                               @                                       @                              @      .@       @                              @                                                      .@       @                                      *@                                               @       @                                       @                                                       @                              6@      D@      H@      $@                      6@     �C@      4@                              ,@     �B@      3@                              $@     �A@      3@                              $@     �@@                                      @      @                                      @      @                                       @      @                                       @                                                      @                                      �?                                              @                                              @      >@                                      @      "@                                      @      �?                                      @                                                      �?                                               @                                              5@                                               @      3@                                              3@                                       @                                      @       @                                      @                                                       @                                       @       @      �?                              @                                              �?       @      �?                                       @                                      �?              �?                                              �?                              �?                                                      �?      <@      $@                              �?      3@      @                                      0@      �?                                      @      �?                                      �?      �?                                      �?                                                      �?                                      @                                              (@                                      �?      @       @                              �?              �?                                              �?                              �?                                                      @      �?                                      @                                                      �?                                      "@      @                                      @                                              @      @                                      @                                                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hKhNhJ	NhG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKՅ�h��B�.         |                    @gy}$x��?�            `u@       i                    �?����?�             k@                           �?����3�?u            `g@                           �?������?            �D@                           �?�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?                           �?��S�ۿ?             >@	       
                     @      �?             0@������������������������       �                     @                           �?�<ݚ�?             "@              #             �?�q�q�?             @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     ,@       :                    @�1�͢S�?Y            @b@       5                    �?z�W�6��?.            @U@                           �?��[����?)            �R@              &             �?�8��8��?             @                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @       *                    �?\��Z���?&            @Q@       #                     @��O�+��?            �E@       "                     �?XB���?             =@              )             �?؇���X�?             @������������������������       �                     @        !       %             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     6@$       '       '             �?؇���X�?	             ,@%       &                    �?      �?              @������������������������       �                     �?������������������������       �                     �?(       )                    �?�8��8��?             (@������������������������       �                     &@������������������������       �                     �?+       ,       %             �?8�Z$���?             :@������������������������       �                     (@-       0                    �?����X�?	             ,@.       /       #             �?      �?             @������������������������       �                      @������������������������       �                      @1       4                    �?z�G�z�?             $@2       3                    �?����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @6       7                    �?���Q��?             $@������������������������       �                     @8       9       !             �?؇���X�?             @������������������������       �                     �?������������������������       �                     @;       ^                    �?0��Jy��?+            �N@<       Y                    �?b�2�tk�?$             K@=       B                    �?8��"���?!            �H@>       A                    �?������?             @?       @       
             �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @C       X                    �?�-�I	p�?             E@D       S                    �?Xތ��?            �D@E       J                    �?     ��?             @@F       G                    �?�nkK�?             7@������������������������       �                     2@H       I                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?K       P       )             �?h/�����?             "@L       M                    �?�$I�$I�?             @������������������������       �                     @N       O       %             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @Q       R                    �?      �?              @������������������������       �                     �?������������������������       �                     �?T       U                    �?X�<ݚ�?             "@������������������������       �                     @V       W                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?Z       ]                    @{�G�z�?             @[       \                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @_       h       $             �?:/����?             @`       e                    �?{�G�z�?             @a       d                    �?�q�q�?             @b       c                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?f       g                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @j       m                    �?���.�?             >@k       l       %             �?8�Z$���?	             *@������������������������       �                     &@������������������������       �                      @n       u                    �?�l� {�?             1@o       t                    @�eP*L��?             &@p       s                     �?r�q��?             @q       r                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @v       y                    @VUUUUU�?             @w       x                     @      �?              @������������������������       �                     �?������������������������       �                     �?z       {                    �?      �?             @������������������������       �                     @������������������������       �                     �?}       �       &             �?�%jj�?O            @_@~       �                    �?R����?4             T@       �                    @��Ņ-]�?'            �M@�       �       '             �?�D�����?             5@�       �       $             �?�8��8��?	             (@�       �                    @      �?              @�       �                    @؇���X�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �       )             �?      �?             @������������������������       �                      @������������������������       �                      @�       �       !             �?�<ݚ�?             "@������������������������       �                     @�       �                     @���Q��?             @������������������������       �                      @������������������������       �                     @�       �                    �?���y4F�?             C@�       �                    �? �Cc}�?             <@������������������������       �        
             3@�       �       #             �?�q�q�?             "@�       �                    @և���X�?             @������������������������       �                     �?�       �       '             �?      �?             @�       �                    �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                    �?      �?             $@�       �                    �?����X�?             @�       �       	             �?r�q��?             @������������������������       �                     @�       �                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �?>4և���?             5@������������������������       �                      @�       �                    �?��uJ���?             3@�       �                    @և���X�?             @������������������������       �                     @������������������������       �                     @�       �                    �?�������?             (@�       �                    �?
ףp=
�?             @�       �                    �?      �?             @������������������������       �                      @�       �                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �?,h��ȓ�?            �F@�       �                    �?Y�����?             &@�       �                    @؇���X�?             @������������������������       �                     @������������������������       �                     �?�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �?�g+��?             A@�       �       !             �?>F?�!��?             5@�       �                    �?<+	���?
             .@�       �                     �?�z�G��?             $@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    @���Q��?             @������������������������       �                      @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    @�8��8��?             @������������������������       �                      @�       �                    @      �?             @������������������������       �                     @������������������������       �                     �?�       �                    @�؉�؉�?             *@�       �                     �?ףp=
�?             $@�       �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�t�bh�h)h,K ��h.��R�(KK�KK��h�B�'        D@      L@     �X@     @T@      H@      3@      :@     �B@      U@      J@      "@      "@      .@      ?@     �R@      J@       @      @      (@      =@                                      $@      �?                                      $@                                                      �?                                       @      <@                                       @      ,@                                              @                                       @      @                                       @      �?                                      �?      �?                                              �?                                      �?                                              �?                                                      @                                              ,@                                      @       @     �R@      J@       @      @      @       @      Q@      (@                      @       @      P@      @                      @      �?       @                                      �?       @                                               @                                      �?                                      @                                                      �?      O@      @                              �?      D@       @                              �?      <@                                      �?      @                                              @                                      �?      �?                                      �?                                                      �?                                              6@                                              (@       @                                      �?      �?                                              �?                                      �?                                              &@      �?                                      &@                                                      �?                                      6@      @                                      (@                                              $@      @                                       @       @                                       @                                                       @                                       @       @                                      @       @                                      @                                                       @                                      @                                              @      @                                      @                                              �?      @                                      �?                                                      @                                      @      D@       @      @                      @      C@      @      @                      @      B@      @      @                              @      �?      @                              @      �?                                      @                                                      �?                                                      @                      @     �@@      @       @                      @     �@@      @       @                      @      ;@       @                              �?      6@                                              2@                                      �?      @                                              @                                      �?                                               @      @       @                              �?      @       @                                      @                                      �?               @                              �?                                                               @                              �?      �?                                      �?                                                      �?                                              @      �?       @                              @                                                      �?       @                                      �?                                                       @                                      �?                               @       @              �?                               @              �?                               @                                                              �?                       @                                               @       @      @                               @       @      �?                              �?       @                                      �?      �?                                              �?                                      �?                                                      �?                                      �?              �?                              �?                                                              �?                                               @              &@      @      "@              �?      @      &@               @                              &@                                                               @                                      @      @              �?      @              @      @                                      @      �?                                      �?      �?                                      �?                                                      �?                                      @                                                      @                                      �?      �?              �?      @              �?      �?                                      �?                                                      �?                                                              �?      @                                              @                                      �?              ,@      3@      ,@      =@     �C@      $@       @       @      @      :@      B@      "@       @       @      @      *@      >@       @       @       @      @      *@                       @              @      @                                       @      @                                      �?      @                                      �?      �?                                      �?                                                      �?                                              @                                      �?                               @               @                               @                                                               @                                       @              @                                              @                               @              @                               @                                                              @                                                      >@       @                                      9@      @                                      3@                                              @      @                                      @      @                                      �?                                              @      @                                       @      @                                       @                                                      @                                      �?                                               @                                              @      @                                       @      @                                      �?      @                                              @                                      �?      �?                                      �?                                                      �?                                      �?                                              @                              �?      *@      @      �?                                       @                              �?      *@      @      �?                              @      @                                      @                                                      @                              �?      "@      �?      �?                      �?       @      �?      �?                               @      �?      �?                               @                                                      �?      �?                                      �?                                                      �?                      �?                                                      @                      (@      1@      "@      @      @      �?      @      �?      @                              @              �?                              @                                                              �?                                      �?      @                                      �?                                                      @                              @      0@      @      @      @      �?      @      @      @       @      @      �?      @      @      @       @                      @      @                                      @      �?                                      @                                                      �?                                              @                                                      @       @                                       @                                              �?       @                                      �?                                                       @                                       @              @      �?                       @                                                              @      �?                                      @                                                      �?      @      "@              �?                              "@              �?                              @              �?                              @                                                              �?                              @                                      @                                        �t�bubhhubh)��}�(hhhhhNhKhKhG        hKhNhJ���%hG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKӅ�h��B(.         �                    @�������?�            `u@       5                    �?BF_�?�            �m@       0                    �?��>4և�?9             U@       #                    �?��y�:�?.            �P@                           �?�[�IJ�?!            �G@������������������������       �                     @                           �?#z�i��?            �D@                           �?r֛w���?             ?@	                           �?8�Z$���?             :@
                           �?�LQ�1	�?             7@                           �?����X�?             @������������������������       �                     �?                            �?r�q��?             @������������������������       �                     @������������������������       �                     �?                           �?      �?	             0@                           �?ףp=
�?             $@������������������������       �                      @              "             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?                           �?z�G�z�?             @              	             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @       "                     �?���Q��?             $@        !                    �?�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @$       -                    @ףp=
�?             4@%       ,                    �?�IєX�?
             1@&       '                    �?�����H�?             "@������������������������       �                     @(       +                    �?�q�q�?             @)       *       )             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @.       /                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?1       2                    �?ҳ�wY;�?             1@������������������������       �                      @3       4                    �?�q�q�?             "@������������������������       �                     @������������������������       �                     @6       y                    �?��p��z�?b             c@7       j                    @6��
J��?<             W@8       Q       #             �?�����2�?0            @Q@9       D                    �?��&��?             9@:       C                    �?�8��8��?             (@;       >                    �?}��7�?             &@<       =                     �?�q�q�?             @������������������������       �                     @������������������������       �                      @?       @       '             �?z�G�z�?             @������������������������       �                     @A       B                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?E       H                    @*D>��?             *@F       G       $             �?      �?             @������������������������       �                     �?������������������������       �                     @I       N                    �?B{	�%��?             "@J       K                     �?r�q��?             @������������������������       �                      @L       M                    @      �?             @������������������������       �                     @������������������������       �                     �?O       P       !             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @R       W                    @�����|�?             F@S       T                    �?$�q-�?             :@������������������������       �                     6@U       V       )             �?      �?             @������������������������       �                      @������������������������       �                      @X       a                    �?)O���?             2@Y       `                    �?      �?              @Z       _                    �?VUUUUU�?             @[       ^                    �?�Q����?             @\       ]                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                      @b       i                    �?p=
ףp�?	             $@c       f                     �?B{	�%��?             "@d       e                    �?؇���X�?             @������������������������       �                     @������������������������       �                     �?g       h                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?k       t       '             �?$G�h��?             7@l       m                    �?     ��?             0@������������������������       �                     @n       s                    @h/�����?             "@o       r                    �?z�G�z�?             @p       q                      @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @u       v       &             �?�$I�$I�?             @������������������������       �                      @w       x       $             �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?z       �                    @ ��i��?&            �N@{       �       
             �?�U��nd�?#             K@|       �                    @�G�z�?             D@}       �       #             �?�<ݚ�?             "@~                           �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �       $             �?�g�y��?             ?@������������������������       �                     5@�       �                    �?ףp=
�?             $@������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �       $             �?և���X�?	             ,@�       �       )             �?����X�?             @�       �                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �?؇���X�?             @������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?����X�?             @������������������������       �                     @������������������������       �                      @�       �                    @��5-p�?=            @Z@�       �                    @㺥��?            �@@�       �                    @0�G�2��?             ;@������������������������       �                     @�       �                    �?���}<S�?             7@������������������������       �                      @������������������������       �                     5@�       �                    �?�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                    �?uk~X��?*             R@�       �       %             �?8�A`���?             I@������������������������       �                     @�       �                    �?��^|��?             G@�       �                    @أp=
��?             D@�       �       
             �?r�q��?             @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �       !             �?H�V�e��?             A@�       �                    �?�IєX�?	             1@������������������������       �                     $@�       �                    �?؇���X�?             @�       �                    @�q�q�?             @������������������������       �                     �?�       �       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    @ҳ�wY;�?
             1@�       �                    �?8�Z$���?             *@�       �                    @�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                     @r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    �?�x?r���?             6@�       �       $             �?p=
ףp�?             $@�       �                    �?      �?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �       	             �?�������?             (@�       �                    �?���Q��?             @������������������������       �                     @������������������������       �                      @�       �                    @����X�?             @������������������������       �                     �?�       �                    �?r�q��?             @�       �                      @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�t�bh�h)h,K ��h.��R�(KK�KK��h�B�'       �B@     �K@     �V@     �U@     �H@      9@     �A@     �K@     @U@     �D@      *@       @     �@@     �I@                                      6@     �F@                                      4@      ;@                                      @                                              ,@      ;@                                       @      7@                                      @      6@                                      @      4@                                       @      @                                      �?                                              �?      @                                              @                                      �?                                              �?      .@                                      �?      "@                                               @                                      �?      �?                                      �?                                                      �?                                              @                                      �?       @                                               @                                      �?                                              @      �?                                      �?      �?                                      �?                                                      �?                                      @                                              @      @                                       @      @                                       @                                                      @                                      @                                               @      2@                                      �?      0@                                      �?       @                                              @                                      �?       @                                      �?      �?                                              �?                                      �?                                                      �?                                               @                                      �?       @                                               @                                      �?                                              &@      @                                       @                                              @      @                                              @                                      @                                               @      @     @U@     �D@      *@       @       @       @      D@      =@      *@      @       @       @     �A@      1@      @      @       @              @      "@       @      @       @              @      �?      �?      @       @              @      �?              @       @                                      @                                              @       @                                                              @      �?                                      @                                              �?      �?                                              �?                                      �?                                                              �?                              @       @      �?      �?                      @      �?                                              �?                                      @                                                      @      �?      �?                              @      �?                                       @                                              @      �?                                      @                                                      �?                                       @              �?                                              �?                               @                               @      <@       @      @      �?               @      8@                                              6@                                       @       @                                       @                                                       @                                              @       @      @      �?                      @      �?      @      �?                      �?      �?      @      �?                              �?      @      �?                              �?              �?                              �?                                                              �?                                      @                              �?                                               @                                              �?      @       @                              �?      @      �?                              �?      @                                              @                                      �?                                                      �?      �?                                              �?                                      �?                                                      �?                              @      (@      @                              �?      &@      @                                      @                                      �?      @      @                              �?      @                                      �?       @                                               @                                      �?                                                       @                                                      @                              @      �?       @                                               @                              @      �?                                      @                                                      �?                               @     �F@      (@               @               @     �F@      @                               @     �B@      �?                               @      @                                       @       @                                               @                                       @                                                      @                                              >@      �?                                      5@                                              "@      �?                                      @                                               @      �?                                       @                                                      �?                                       @      @                                       @      @                                       @      �?                                       @                                                      �?                                              @                                      @      �?                                      @                                              �?      �?                                              �?                                      �?                                                      @               @                              @                                                               @       @              @     �F@      B@      1@                      @      5@      @      @                      @      5@       @                              @                                                      5@       @                                               @                                      5@                                                       @      @                                              @                                       @               @              �?      8@      @@      *@                      �?      ,@      <@      @                              @                                      �?      $@      <@      @                      �?      @      ;@      @                      �?      @                                              @                                      �?       @                                               @                                      �?                                                              ;@      @                                      0@      �?                                      $@                                              @      �?                                       @      �?                                      �?                                              �?      �?                                      �?                                                      �?                                      @                                              &@      @                                      &@       @                                      $@      �?                                      $@                                                      �?                                      �?      �?                                      �?                                                      �?                                              @                              @      �?                                      @                                                      �?               @                      $@      @      @                              @       @      �?                              �?       @      �?                              �?              �?                                              �?                              �?                                                       @                                      @                       @                      @       @      @       @                      @                                              @                       @                                                                               @      @                                      �?                                              �?      @                                      �?       @                                      �?                                                       @                                              @�t�bubhhubh)��}�(hhhhhNhKhKhG        hKhNhJs-hG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK���h��B�(         ,                    �?�zz*l��?�            `u@                           �?l��[B��?<            �U@                           �?ܷ��?��?             =@              
             �? ��WV�?             :@������������������������       �                     7@                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @	       
                     �?�q�q�?             @������������������������       �                      @������������������������       �                     �?       '                    �?�c�Α�?+             M@       "                    �?�㙢�c�?%             G@                           �?�ݜ�?            �C@������������������������       �                     �?                            @�KM�]�?             C@                           �? 7���B�?             ;@������������������������       �                     6@                           �?z�G�z�?             @                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @       !                    �?���!pc�?	             &@              #             �?      �?             @                           �?      �?             @                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?                            �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @#       &                     �?և���X�?             @$       %                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @(       +                     @�q�q�?             (@)       *                    �?z�G�z�?             $@������������������������       �                      @������������������������       �                      @������������������������       �                      @-       �                    @�=����?�            �o@.       ]       %             �?>wOE=l�?�            �k@/       V                    �?�w#�z&�?5            @U@0       M                    @Z2���h�?/             S@1       L       	             �?��9�D�?$            �L@2       9                     �?J�$I�$�?#             L@3       6                    @������?             ,@4       5                    �?z�G�z�?             $@������������������������       �                      @������������������������       �                      @7       8                    �?      �?             @������������������������       �                     @������������������������       �                     �?:       K                    �?����S�?             E@;       J                    �?أp=
��?             D@<       =                    �?dG�+�?             ?@������������������������       �                     �?>       E                    �?�h$���?             >@?       D                    �?���N8�?             5@@       C                    @ףp=
�?             $@A       B       "             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     &@F       G                    �?�<ݚ�?             "@������������������������       �                     @H       I       !             �?�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     "@������������������������       �                      @������������������������       �                     �?N       U                    @0\�Uo��?             3@O       R                    �?��1G���?             *@P       Q                    �?���Q��?             @������������������������       �                      @������������������������       �                     @S       T                    �?      �?              @������������������������       �                      @������������������������       �                     @������������������������       �                     @W       Z                    �?��E���?             "@X       Y                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?[       \                     �?�q�q�?             @������������������������       �                      @������������������������       �                     �?^       _                    @�9�?Q            �`@������������������������       �        
             0@`       �                    �?���S���?G            �]@a       �                    �? �\�Y��?@            �Z@b       q                    �?���W��?3            @T@c       h                    �?x�"w���?             3@d       g                    @0�����?             @e       f                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?i       n                    �?9��8���?             (@j       k                    �?0�����?             @������������������������       �                     �?l       m                    �?r�q��?             @������������������������       �                     �?������������������������       �                     @o       p       !             �?���Q��?             @������������������������       �                     @������������������������       �                      @r       �                    �?0LbOV��?&             O@s       |                     �?<73V�=�?#            �L@t       w                    �?X�Cc�?             ,@u       v                    �?      �?             @������������������������       �                     �?������������������������       �                     @x       {                    @z�G�z�?             $@y       z                    @�����H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �                     �?}       �                    �?���*�?            �E@~       �                    @���y4F�?             C@       �       "             �?\-��p�?             =@�       �                    @���y4F�?             3@������������������������       �                     *@�       �       $             �?�q�q�?             @�       �                    �?      �?             @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@�       �       !             �?X�<ݚ�?             "@�       �                    �?�q�q�?             @�       �                    @�q�q�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �?{�G�z�?             @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    @��%��?             :@�       �                    �?      �?             8@�       �                    @�nkK�?             7@�       �                     �?؇���X�?             @�       �                    @      �?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     0@������������������������       �                     �?������������������������       �                      @�       �       "             �?r�q��?             (@�       �                    �?���(\��?             $@�       �                    �?X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                    @�E����?            �A@�       �                    @؇���X�?             5@�       �                     @ףp=
�?             4@������������������������       �                     0@�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?�       �                    �?�X�C�?
             ,@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    @�eP*L��?             &@������������������������       �                     @������������������������       �                     @�t�bh�h)h,K ��h.��R�(KK�KK��h�B#       �E@     �K@      T@     �W@     �I@      2@      E@     �F@                                      :@      @                                      9@      �?                                      7@                                               @      �?                                              �?                                       @                                              �?       @                                               @                                      �?                                              0@      E@                                       @      C@                                      @      A@                                      �?                                              @      A@                                      �?      :@                                              6@                                      �?      @                                      �?       @                                      �?                                                       @                                               @                                      @       @                                      @      @                                       @       @                                       @      �?                                              �?                                       @                                                      �?                                      �?      �?                                      �?                                                      �?                                              @                                      @      @                                      @      �?                                              �?                                      @                                                      @                                       @      @                                       @       @                                       @                                                       @                                               @                                      �?      $@      T@     �W@     �I@      2@      �?      $@      T@     @W@      <@       @      �?      @     �I@      6@      @      @      �?      @      I@      1@       @       @      �?      @      F@       @                      �?      @      F@      @                              @       @      @                               @       @                                       @                                                       @                                      �?              @                                              @                              �?                                      �?      �?      B@      @                      �?      �?      B@       @                      �?      �?      ;@       @                      �?                                                      �?      ;@       @                              �?      4@                                      �?      "@                                      �?       @                                               @                                      �?                                                      @                                              &@                                              @       @                                      @                                              @       @                                      @                                                       @                                      "@                                                       @                                              �?                                      @      "@       @       @                      @      @       @       @                              @       @                                               @                                      @                                      @                       @                                               @                      @                                                      @                                      �?      @       @      �?                      �?      @                                              @                                      �?                                                               @      �?                                       @                                                      �?              @      =@     �Q@      8@      @                      0@                                      @      *@     �Q@      8@      @               @       @     @Q@      7@      @               @      @     �G@      5@      @                      @      @      @      @                      �?      @              �?                      �?      @                                              @                                      �?                                                                      �?                      @              @      @                      @              �?      �?                                              �?                      @              �?                                              �?                              @                                                              @       @                                      @                                                       @               @      �?      E@      1@                       @      �?     �B@      1@                                      @      "@                                      @      �?                                              �?                                      @                                               @       @                                      �?       @                                      �?                                                       @                                      �?                               @      �?      @@       @                                      >@       @                                      9@      @                                      .@      @                                      *@                                               @      @                                       @       @                                       @      �?                                              �?                                       @                                                      �?                                               @                                      $@                                              @      @                                       @      @                                       @      �?                                      �?      �?                                      �?                                                      �?                                      �?                                                      @                                      @                               @      �?       @                               @      �?                                       @                                                      �?                                                       @                                              @                                      �?      6@       @      �?                      �?      6@              �?                      �?      6@                                      �?      @                                      �?      @                                      �?      �?                                              �?                                      �?                                                       @                                              @                                              0@                                                              �?                                       @                      @      @       @      �?                      @      @              �?                      @      @                                              @                                      @                                                                      �?                                       @                                               @      7@      $@                                      2@      @                                      2@       @                                      0@                                               @       @                                       @                                                       @                                              �?                               @      @      @                               @              �?                                              �?                               @                                                      @      @                                      @                                                      @�t�bub�?     hhubh)��}�(hhhhhNhKhKhG        hKhNhJ�E^hG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKǅ�h��B�+         ~                    @��Hs��?�            `u@       9       &             �?�hw�G�?�            �l@       8                    @�d�Y��?5            �U@       /                    @k�=F?��?4             U@       .                    �?*�	�3�?+            @Q@              #             �?{�����?(            @P@                           �?&���^B�?             2@                           �?H�7�&��?             .@	                           �?{�G�z�?             @
                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     $@                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?       !       
             �?�rCzA��?            �G@                           �?VUUUUU�?             8@                           @���Q��?             $@������������������������       �                     @                           �?؇���X�?             @������������������������       �                     @                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?                            �?0�����?             ,@                           �?r�q��?             (@                           �?�<ݚ�?             "@������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                      @"       )                    �?H��	,U�?             7@#       $                    @>;n,��?             &@������������������������       �                     @%       (                     �?0�����?             @&       '                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @*       +                    �?r�q��?             (@������������������������       �                      @,       -                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @0       1                     @��S���?	             .@������������������������       �                     @2       3       
             �?z�G�z�?             $@������������������������       �                     �?4       5                    �?�����H�?             "@������������������������       �                     @6       7                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @:       I                     �?�qM{���?Q            �a@;       @       )             �?hha�H��?             =@<       ?                    �?���Q��?             .@=       >                    �?@4և���?             ,@������������������������       �                     *@������������������������       �                     �?������������������������       �                     �?A       H                    �?�$I�$I�?             ,@B       G                     �?      �?             (@C       D                    @z�G�z�?             $@������������������������       �                     @E       F                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                      @J       _                    �?�Z�?D            @\@K       L                    �?Fmq��?"            �J@������������������������       �                     *@M       ^       !             �?z�G�z�?             D@N       Y                    �?�	j*D�?             :@O       X                    �?���y4F�?             3@P       U       
             �?�t����?             1@Q       R                    �?��S�ۿ?	             .@������������������������       �                      @S       T                     �?؇���X�?             @������������������������       �                     @������������������������       �                     �?V       W       '             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @Z       ]                    �?և���X�?             @[       \                    �?�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �        	             ,@`       g                    �?�������?"             N@a       f                    �?
ףp=
�?             $@b       e                    �?VUUUUU�?             "@c       d                    �?      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     �?h       y                    �?Ǻ���?             I@i       x       (             �?h\�A�
�?            �F@j       u                    �?��O�+��?            �E@k       n       "             �?x1z�?�?            �C@l       m                    @�g�y��?             ?@������������������������       �                     >@������������������������       �                     �?o       t                    �?      �?              @p       q                    �?z�G�z�?             @������������������������       �                      @r       s                    @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @v       w                    @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @z       {                     @���Q��?             @������������������������       �                      @|       }       #             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?       �                    @�1�g
�?M            @\@�       �       %             �?��_�}�?-             Q@�       �                    �?6������?            �C@�       �                    �?�z�G��?             4@�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @�       �                    �?      �?             0@�       �       )             �?z�G�z�?
             .@������������������������       �                     @�       �       
             �?      �?              @������������������������       �                     @�       �       	             �?���Q��?             @������������������������       �                     �?�       �                     �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?�       �                    �?��|���?             3@�       �                    �?ƒ_,���?
             .@�       �                    @/y0��k�?	             *@�       �                    �?�z�G��?             $@������������������������       �                     @�       �                    �?���Q��?             @������������������������       �                     �?�       �                      @      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �?�8���?             =@�       �                    �?�eP*L��?             6@������������������������       �                     �?�       �                     @�E�_���?             5@�       �                    �?VUUUUU�?             @�       �       #             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �        
             2@�       �       )             �?և���X�?             @������������������������       �                      @�       �                    �?z�G�z�?             @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �       %             �?������?             �F@�       �       
             �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?>��C��?            �E@�       �                    �?ףp=
�?             4@�       �                    �?�X�<ݺ?             2@������������������������       �        	             ,@�       �       "             �?      �?             @������������������������       �                     @������������������������       �                     �?�       �       
             �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �       $             �?�LQ�1	�?             7@�       �                    @     ��?
             0@������������������������       �                     *@������������������������       �                     @�       �                    @����X�?             @������������������������       �                     �?�       �                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?�t�bh�h)h,K ��h.��R�(KK�KK��h�BP%        F@     �N@     �T@     �S@      K@      5@     �B@      G@     @Q@      H@      3@      $@               @      4@      D@      2@      @               @      4@      D@      .@      @               @      4@      D@      @                       @      4@      B@      @                              �?      *@      @                              �?      (@       @                              �?       @       @                              �?               @                              �?                                                               @                                       @                                              $@                                              �?       @                                               @                                      �?                               @      3@      7@      @                       @      ,@       @                                      @      @                                      @                                              �?      @                                              @                                      �?       @                                               @                                      �?                                       @      $@       @                                      $@       @                                      @       @                                      @                                                       @                                      @                                       @                                                      @      .@      @                              @      @      �?                              @                                              �?      @      �?                              �?              �?                              �?                                                              �?                                      @                                              $@       @                                       @                                               @       @                                       @                                                       @                                      @                                                       @      @                                              @                                       @       @                                              �?                                       @      �?                                      @                                              @      �?                                      @                                                      �?                                      @             �B@      F@     �H@       @      �?      @      *@      "@      @      @                      *@      �?      �?                              *@      �?                                      *@                                                      �?                                                      �?                                       @       @      @                               @       @       @                               @               @                              @                                               @               @                                               @                               @                                                       @                                                       @                      8@     �A@      G@      @      �?      @      5@      @@                                      *@                                               @      @@                                       @      2@                                      @      .@                                       @      .@                                      �?      ,@                                               @                                      �?      @                                              @                                      �?                                              �?      �?                                      �?                                                      �?                                       @                                              @      @                                      @       @                                      @                                                       @                                              �?                                              ,@                                      @      @      G@      @      �?      @      @              @              �?      @      @              @                      @      @                                      @      @                                                                                      @                      @                                                              �?                      @     �E@      @                              @      D@       @                              �?      D@       @                              �?     �B@      �?                                      >@      �?                                      >@                                                      �?                              �?      @                                      �?      @                                               @                                      �?       @                                      �?                                                       @                                              @                                              @      �?                                      @                                                      �?                               @                                                      @       @                                       @                                              �?       @                                               @                                      �?                              @      .@      ,@      ?@     �A@      &@      @      .@      ,@      >@       @              @      ,@      "@       @       @              @      ,@                                       @       @                                               @                                       @                                              @      (@                                      @      (@                                              @                                      @      @                                              @                                      @       @                                      �?                                               @       @                                       @                                                       @                                      �?                                                              "@       @       @                              @       @       @                              @       @       @                              @      @                                              @                                      @       @                                              �?                                      @      �?                                              �?                                      @                                                      �?       @                                               @                                      �?                                       @                                              @                              �?      �?      @      6@                      �?      �?      �?      3@                              �?                                      �?              �?      3@                      �?              �?      �?                      �?              �?                              �?                                                              �?                                                      �?                                              2@                                      @      @                                               @                                      @      �?                                       @      �?                                              �?                                       @                                               @                                                      �?     �@@      &@                              �?              �?                                              �?                              �?                                                     �@@      $@                                      2@       @                                      1@      �?                                      ,@                                              @      �?                                      @                                                      �?                                      �?      �?                                              �?                                      �?                                              .@       @                                      *@      @                                      *@                                                      @                                       @      @                                      �?                                              �?      @                                              @                                      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hKhNhJ�&UhG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKم�h��Bx/         �                    @�(���?�            `u@       E       &             �?�)��?�            �m@       8       "             �?����Mb�?A             Y@                           @S��-fe�?4            �S@                           �?��i~��?            �B@                           @:/����?             5@       
                    @�IєX�?             1@       	                    �?؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     $@              !             �?      �?             @                            �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?                           �?     @�?	             0@                           �?�q�q�?             "@                           �?؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @                           @և���X�?             @������������������������       �                     @                           �?      �?             @������������������������       �                     @������������������������       �                     �?       +                    @��>4և�?             E@       &                    �?Ra���i�?             6@       %       
             �?������?
             1@                             @      �?              @������������������������       �                     @!       $                    �?z�G�z�?             @"       #                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@'       (       '             �?{�G�z�?             @������������������������       �                     �?)       *                     �?      �?             @������������������������       �                      @������������������������       �                      @,       5                    �?���(\��?             4@-       .                    �?     @�?
             0@������������������������       �                     @/       0                    �?޾�z�<�?	             *@������������������������       �                     "@1       2       )             �?      �?             @������������������������       �                      @3       4                     @      �?              @������������������������       �                     �?������������������������       �                     �?6       7                     �?      �?             @������������������������       �                     @������������������������       �                     �?9       D                    @�G��l��?             5@:       =       
             �?9��8���?	             (@;       <                    �?���Q��?             @������������������������       �                      @������������������������       �                     @>       ?                    @�$I�$I�?             @������������������������       �                      @@       C                     �?z�G�z�?             @A       B                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     "@F       �                    �?Z J�P�?[            `a@G       x                    @���-s��?U            ``@H       e                    �?L�y�=�?7            @U@I       L                    �?��Q:��?(            �M@J       K                    �?�8��8��?	             (@������������������������       �                     &@������������������������       �                     �?M       P                    �?��|�5��?            �G@N       O                    �?��S�ۿ?	             .@������������������������       �                     ,@������������������������       �                     �?Q       \                    �?     ��?             @@R       W       #             �?և���X�?	             ,@S       V       $             �?r�q��?             @T       U                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @X       [                    �?      �?              @Y       Z                    �?����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?]       ^       )             �?�����H�?             2@������������������������       �                     $@_       d                    �?      �?              @`       a                    �?؇���X�?             @������������������������       �                     @b       c                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?f       q                    �?Z�K8�?             :@g       l                    �?r�q��?             (@h       k                     �?      �?             @i       j       "             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @m       p                    �?      �?              @n       o       !             �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @r       s                     @@4և���?             ,@������������������������       �                     @t       u                    @؇���X�?             @������������������������       �                     @v       w                    @      �?             @������������������������       �                     �?������������������������       �                     @y       ~                     �?~<SvL�?             G@z       }                    �?      �?              @{       |                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @       �                     @Vo����?             C@�       �                    �?��%��?             :@�       �                    �?�����?             5@������������������������       �                     (@�       �                    �?�<ݚ�?             "@������������������������       �                     @�       �                    �?      �?             @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                     �?�Q����?             @�       �                     @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �?9��8���?	             (@�       �                    �?z�G�z�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �       #             �?և���X�?             @������������������������       �                     @������������������������       �                     @�       �       !             �?      �?              @�       �                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                     @      �?              @������������������������       �                     �?������������������������       �                     �?�       �       	             �?;p����?E            �Y@�       �                    @������?4            �S@�       �                     @�Xi�|.�?%            �L@�       �                    @����?             7@�       �       !             �?�q�q�?	             (@�       �       )             �?r�q��?             @�       �       &             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                      @�       �       '             �?      �?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    @���!pc�?             &@�       �                    �?      �?             @�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �?hJ,���?             A@�       �                    �?dG�+�?             ?@�       �                    �?P���Q�?             4@������������������������       �                     3@������������������������       �                     �?�       �                    �?j�V���?             &@�       �                    @�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                    @�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?"pc�
�?             6@�       �                    @���Q��?             @������������������������       �                     @������������������������       �                      @�       �                    �?�t����?             1@�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �        	             *@�       �                    @9��8���?             8@�       �       %             �?������?
             ,@�       �       #             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?j�V���?             &@�       �                    @z�G�z�?             $@�       �                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     $@�t�bh�h)h,K ��h.��R�(KK�KK��h�B�(        C@      P@     @S@     �S@     �K@      =@     �B@      N@     @R@      D@      1@      (@      @       @      =@     �@@      0@      &@      @       @      =@      3@      (@       @      @       @      8@       @                               @      1@       @                              �?      0@                                      �?      @                                              @                                      �?                                                      $@                                      �?      �?       @                                      �?       @                                      �?                                                       @                              �?                                      @      @      @                                      @      @                                      @      �?                                      @                                                      �?                                               @                              @              @                                              @                              @              �?                              @                                                              �?                                              @      1@      (@       @                      @      .@       @                              @      *@                                      @      @                                              @                                      @      �?                                      @      �?                                      @                                                      �?                                      �?                                                      "@                                      �?       @       @                              �?                                                       @       @                                       @                                                       @                                       @      $@       @                              �?      $@      @                                              @                              �?      $@       @                                      "@                                      �?      �?       @                                               @                              �?      �?                                      �?                                                      �?                                      �?              @                                              @                              �?                                              ,@      @      @                              @      @      @                              @               @                                               @                              @                                               @      @      �?                               @                                                      @      �?                                      �?      �?                                              �?                                      �?                                              @                                      "@                      A@      J@      F@      @      �?      �?      =@      J@     �E@      @              �?      8@     �E@      .@       @              �?      6@     �B@                                      &@      �?                                      &@                                                      �?                                      &@      B@                                      �?      ,@                                              ,@                                      �?                                              $@      6@                                       @      @                                      @      �?                                      �?      �?                                      �?                                                      �?                                      @                                              @      @                                       @      @                                       @                                                      @                                      �?                                               @      0@                                              $@                                       @      @                                      �?      @                                              @                                      �?      �?                                              �?                                      �?                                              �?                                               @      @      .@       @              �?       @      @       @      �?              �?                       @      �?              �?                              �?              �?                              �?                                                              �?                       @                               @      @                                       @      @                                       @                                                      @                                              @                                                      *@      �?                                      @                                              @      �?                                      @                                              @      �?                                              �?                                      @                              @      "@      <@      @                      @      @      �?                                      @      �?                                      @                                                      �?                              @                                               @      @      ;@      @                       @      �?      6@      �?                       @              3@                                              (@                               @              @                                              @                               @               @                               @              �?                               @                                                              �?                                              �?                                      �?      @      �?                              �?              �?                              �?                                                              �?                                      @                                      @      @      @                              @      �?                                      �?      �?                                              �?                                      �?                                              @                                                      @      @                                              @                                      @                              @              �?      �?      �?              @                      �?                      @                                                                      �?                                      �?              �?                                              �?                              �?                              �?      @      @     �C@      C@      1@              @      @     �A@      >@      @              @      @     �A@      (@      @               @       @      @      "@      @               @       @      @      �?                              �?      @                                      �?       @                                               @                                      �?                                                      @                               @      �?       @      �?                                       @                               @      �?              �?                              �?              �?                              �?                                                              �?                       @                                                                       @      @                                      @      @                                      @      �?                                      @                                                      �?                                               @                                      @                       @      �?      <@      @                       @      �?      ;@      �?                              �?      3@                                              3@                                      �?                                       @               @      �?                                       @      �?                                       @                                                      �?                       @                                                              �?       @                                      �?                                                       @                                              2@      @                                      @       @                                      @                                                       @                                      .@       @                                       @       @                                               @                                       @                                              *@              �?              �?      @       @      $@      �?              �?      @       @                              �?       @                                      �?                                                       @                      �?                       @       @                                       @       @                                       @      �?                                       @                                                      �?                                              @              �?                                                                                      $@�t�bubhhubh)��}�(hhhhhNhKhKhG        hKhNhJ�uhG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKׅ�h��B/         Z                    �?���e�?�            `u@                           �?t��k��?[            �`@                           �?|��?���?$             K@                            @�����?             C@                            �?���Q��?             9@                           �?և���X�?             ,@������������������������       �                     @������������������������       �                      @	                           �?"pc�
�?             &@
                           �?ףp=
�?             $@������������������������       �                     @                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?                           �?8�Z$���?             *@              '             �?      �?              @������������������������       �                     �?������������������������       �                     �?                           @�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?                           �?      �?             0@������������������������       �                     "@                           @����X�?             @                           �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @       Q                    �?>
ףp}�?7             T@       D                    �?��:�
�?(            �M@        9                    �?f+��?            �E@!       8                    @      �?             @@"       +                    @� ��w��?             =@#       *                    @���Q��?             .@$       %                    �?@4և���?
             ,@������������������������       �                     "@&       )                    �?z�G�z�?             @'       (       $             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     �?,       3                    �?����>4�?
             ,@-       0       %             �?�n���?             "@.       /       (             �?      �?             @������������������������       �                      @������������������������       �                      @1       2       '             �?���Q��?             @������������������������       �                      @������������������������       �                     @4       5                    @���Q��?             @������������������������       �                      @6       7                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @:       A                    �?��!pc�?             &@;       @                     @      �?              @<       =                    �?؇���X�?             @������������������������       �                     @>       ?                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?B       C                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @E       P                    �?      �?
             0@F       G                    �?�8��8��?	             (@������������������������       �                     @H       O                     @9��8���?             @I       N                      @      �?             @J       M       !             �?VUUUUU�?             @K       L                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @R       S                    @L�p.0�?             5@������������������������       �                     1@T       Y                    �?      �?             @U       V       $             �?�q�q�?             @������������������������       �                     �?W       X                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?[       �       &             �?��s�.�?{             j@\       k                    �?�*��y�?E            �]@]       h       (             �?�^)��?             9@^       a                    @�X����?             6@_       `                    �?$�q-�?	             *@������������������������       �                     �?������������������������       �                     (@b       g                    �?�n���?             "@c       f       $             �?և���X�?             @d       e                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                      @i       j                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?l       �                    @�DO���?5            �W@m       p                    �?1EYm��?            �I@n       o                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?q       �       )             �?d-<�Z�?            �F@r                            �?�(\����?             4@s       |                    �?�Kh/���?             2@t       u       
             �?/y0��k�?	             *@������������������������       �                     �?v       {                    �?      �?             (@w       z                    @j�V���?             &@x       y       !             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?}       ~                    �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @�       �                    �?���H�?             9@�       �                    @p=
ףp�?
             4@������������������������       �                      @�       �                    @�������?             (@������������������������       �                      @�       �                    �?      �?             @�       �                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �       '             �?��^��?            �E@�       �                    @�\��N��?             3@�       �                    @؇���X�?             @������������������������       �                     @������������������������       �                     �?�       �       !             �?      �?             (@�       �                    �?���!pc�?             &@������������������������       �                     �?�       �                     �?�z�G��?             $@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                    �?�q�q�?             8@�       �       $             �?�d�����?	             3@�       �                    �?�X�<ݺ?             2@������������������������       �                     @�       �                    �?$�q-�?             *@������������������������       �                     @�       �                    �?      �?              @�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                    @���Q��?             @������������������������       �                     @������������������������       �                      @�       �                    �?Y����?6            @V@�       �                    �?�9����?,            �R@�       �       )             �?և���X�?             5@�       �                    �?X�Cc�?
             ,@�       �                    �?�q�q�?             @������������������������       �                     �?�       �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    @      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    �?�Wv���?             K@�       �                    �?�L���o�?            �D@�       �                    @B+K&:~�?             3@�       �       $             �?������?
             1@�       �                    �?����X�?             ,@�       �                    �?���Q��?             $@�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �                    �?�X����?             6@�       �                    �?r�q��?	             2@�       �                     �?      �?             0@������������������������       �                     .@������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �?$�q-�?             *@������������������������       �                     "@�       �       (             �?      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �?�X�C�?
             ,@�       �                    �?      �?	             (@������������������������       �                     @�       �                    @      �?              @�       �                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�t�bh�h)h,K ��h.��R�(KK�KK��h�BP(        G@      H@     �U@      S@      N@      :@      >@      >@     �@@      2@      *@      $@      <@      :@                                      :@      (@                                      .@      $@                                      @       @                                      @                                                       @                                      "@       @                                      "@      �?                                      @                                               @      �?                                              �?                                       @                                                      �?                                      &@       @                                      �?      �?                                      �?                                                      �?                                      $@      �?                                      $@                                                      �?                                       @      ,@                                              "@                                       @      @                                       @       @                                               @                                       @                                                      @                                       @      @     �@@      2@      *@      $@       @      @      0@      0@      (@      "@              @      0@      "@      &@      @              �?      .@      @      @      @              �?      .@      @       @      @              �?      *@      �?                              �?      *@                                              "@                                      �?      @                                      �?       @                                      �?                                                       @                                               @                                                      �?                                       @      @       @      @                       @      @              @                       @                       @                       @                                                                       @                              @               @                                               @                              @                                              @       @                                       @                                              �?       @                                               @                                      �?                                                      @                       @      �?       @      @                                       @      @                                      �?      @                                              @                                      �?      �?                                      �?                                                      �?                                      �?                               @      �?                                              �?                                       @                                       @      �?              @      �?      @       @      �?              @      �?      �?                              @                       @      �?              �?      �?      �?              �?              �?      �?      �?              �?              �?      �?                                      �?      �?                                      �?                                                      �?                      �?                                                                              �?       @                                                                                      @                      1@       @      �?      �?                      1@                                                       @      �?      �?                               @      �?                                      �?                                              �?      �?                                      �?                                                      �?                                                      �?      0@      2@     �J@      M@     �G@      0@                      5@     �B@     �G@      ,@                      @      0@      @                              @      0@      @                              �?      (@                                      �?                                                      (@                                       @      @      @                                      @      @                                      @      �?                                      @                                                      �?                                               @                               @                                               @              �?                               @                                                              �?                              0@      5@     �E@      ,@                      0@      4@      ,@      �?                                      @      �?                                      @                                                      �?                      0@      4@      "@                              @      @       @                              @      @       @                               @      @       @                                      �?                                       @       @       @                               @      �?       @                               @      �?                                       @                                                      �?                                                       @                                      �?                                      @       @                                      @                                                       @                                       @                                              "@      .@      �?                              "@      $@      �?                               @                                              �?      $@      �?                                       @                                      �?       @      �?                                       @      �?                                       @                                                      �?                              �?                                                      @                                              �?      =@      *@                                      "@      $@                                      @      �?                                      @                                                      �?                                      @      "@                                      @       @                                              �?                                      @      @                                      @      �?                                      @                                                      �?                                              @                                              �?                              �?      4@      @                              �?      1@      �?                                      1@      �?                                      @                                              (@      �?                                      @                                              @      �?                                      @      �?                                      @                                                      �?                                      @                                      �?                                                      @       @                                      @                                                       @      0@      2@      @@      5@               @      "@      *@      @@      3@               @      "@      (@                                      "@      @                                       @      @                                      �?                                              �?      @                                              @                                      �?                                              @      �?                                      @                                                      �?                                              @                                              �?      @@      3@               @                      4@      3@               @                      *@      @               @                      *@      @                                      $@      @                                      @      @                                      �?      @                                      �?                                                      @                                      @                                              @                                              @                                                                       @                      @      .@                                      @      .@                                      �?      .@                                              .@                                      �?                                               @                                              @                                      �?      (@                                              "@                                      �?      @                                              @                                      �?                                      @      @               @                      @      @               @                      @                                              �?      @               @                      �?      @                                              @                                      �?                                                                       @                       @                                        �t�bub��      hhubh)��}�(hhhhhNhKhKhG        hKhNhJ�G5GhG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKh��BH4         �                    �?F�f%��?�            `u@       }                    �?�/�\m;�?�             p@       6       &             �?ܰe?��?x            �g@       %                    @ 2�P���?/            @S@                           �?_�#���?              K@                           @/�����?             <@                            �?�"�O�|�?             1@       	                    �?{�G�z�?             @������������������������       �                      @
              )             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     (@                           �?���!pc�?             &@������������������������       �                     @                           �?���Q��?             @������������������������       �                     @������������������������       �                      @       "                     @g\�5�?             :@                           �?     ��?
             0@                           �?��8��8�?             (@                           �?      �?              @                           @      �?             @              '             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @                           �?      �?             @������������������������       �                     @������������������������       �                     �?        !       $             �?      �?             @������������������������       �                     @������������������������       �                     �?#       $                     @ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@&       /                    �?
;&����?             7@'       ,                    @>;n,��?             &@(       +                     �?r�q��?             @)       *       #             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @-       .                     @z�G�z�?             @������������������������       �                     @������������������������       �                     �?0       1       )             �?�������?             (@������������������������       �                      @2       5                    �?      �?             @3       4                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?7       z       	             �?�"QQ(��?I            @\@8       g                     �?&K:�m��?F             [@9       <                    �?��87d�?2            @S@:       ;                    @r�q��?             @������������������������       �                     @������������������������       �                     �?=       P                    �?.c!�?-            �Q@>       K                    �?���Q��?             >@?       J                    @�GN�z�?             6@@       I                    �?�E��ӭ�?             2@A       B                    �?     ��?             0@������������������������       �                      @C       H       #             �?@4և���?             ,@D       E                    �?z�G�z�?             @������������������������       �                     @F       G       $             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@������������������������       �                      @������������������������       �                     @L       O                    �?      �?              @M       N       '             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @Q       `                    �?��d;�w�?            �D@R       [                    @z5�h$�?             >@S       Z                    @      �?             4@T       U                     @      �?
             0@������������������������       �                     $@V       W                    �?r�q��?             @������������������������       �                     @X       Y       "             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @\       ]                    �?H�z�G�?             $@������������������������       �                     @^       _                    �?      �?             @������������������������       �                     @������������������������       �                     �?a       f                     @�C��2(�?             &@b       c                    �?      �?             @������������������������       �                      @d       e       "             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @h       m                    �?~eC����?             ?@i       j                    �?�C��2(�?             &@������������������������       �                     @k       l                    �?      �?             @������������������������       �                     �?������������������������       �                     @n       y       )             �?H�z�G�?             4@o       x                    �?8�Z$���?	             *@p       s                    @j�V���?             &@q       r       
             �?      �?              @������������������������       �                     �?������������������������       �                     �?t       w                    �?�����H�?             "@u       v                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @{       |                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?~       �                    �?�G�V�e�?1             Q@       �       "             �?��k���?             F@�       �       &             �?�Q����?             D@�       �                     @�E]t��?             6@�       �                    �?I�$I�$�?             ,@�       �                    �?�<ݚ�?             "@�       �                    �?      �?              @�       �                    �?      �?             @�       �                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                    �?{�G�z�?             @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                      @�       �       )             �?h/�����?             2@�       �                    @��ˠ�?	             &@������������������������       �                     @�       �                    �?      �?              @�       �       !             �?0�����?             @�       �                     @VUUUUU�?             @������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �       !             �?����X�?             @������������������������       �                     @�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @�       �                    �?      �?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �       "             �?�q�q�?             8@�       �                    �?F]t�E�?             6@�       �                    �?�l� {�?             1@�       �                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    @������?	             &@�       �       $             �?������?             @�       �                    @�Q����?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                     �?      �?             @������������������������       �                     �?������������������������       �                     @�       �       (             �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @�       �                    @	p��&%�?1             U@�       �                     �?pX���o�?"            �K@�       �                     @���O]�?            �B@�       �                    @�u]�u]�?             5@�       �                    �?�8��8��?             (@�       �                    @X�<ݚ�?             "@������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    @VUUUUU�?             "@�       �                    �?�Q����?             @������������������������       �                     �?�       �       
             �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    @      �?             0@�       �                    �?VUUUUU�?             @�       �       "             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                    �?$�q-�?             *@������������������������       �                     �?������������������������       �                     (@�       �                    @n�����?	             2@�       �       &             �?�2�tk~�?             "@�       �                    @�q�q�?             @������������������������       �                      @�       �       #             �?      �?             @������������������������       �                     �?�       �                    @�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �       "             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                     @�<ݚ�?             "@������������������������       �                      @������������������������       �                     @�       �                    @J�8���?             =@�       �                    @��<b���?             7@������������������������       �        
             2@������������������������       �                     @�       �       
             �?r�q��?             @������������������������       �                     �?������������������������       �                     @�t�bh�h)h,K ��h.��R�(KK�KK��h�B�,        C@      J@     �V@     �R@     @P@      6@      A@     �H@      T@      K@      A@      @      ?@     �@@     �P@      E@      0@       @       @      @      6@      ?@      .@       @       @      @      6@      9@                               @      1@      "@                               @      ,@      �?                               @       @      �?                               @                                                       @      �?                                       @                                                      �?                                      (@                                              @       @                                              @                                      @       @                                      @                                                       @                       @      @      @      0@                      �?      @      @      @                      �?              @      @                                      @      @                                      �?      @                                      �?      �?                                              �?                                      �?                                                       @                                      @                              �?                      @                                              @                      �?                                                      @              �?                              @                                                              �?                      �?                      "@                      �?                                                                      "@                                              @      .@       @                              @      @      �?                              �?      @                                      �?      �?                                              �?                                      �?                                                      @                                      @              �?                              @                                                              �?                              �?      $@      �?                                       @                                      �?       @      �?                                       @      �?                                       @                                                      �?                              �?                      =@      <@      F@      &@      �?              <@      8@      F@      &@      �?              1@      4@      <@      &@      �?              @      �?                                      @                                                      �?                                      (@      3@      <@      &@      �?              (@      2@                                      @      1@                                      @      *@                                      @      *@                                       @                                              �?      *@                                      �?      @                                              @                                      �?      �?                                      �?                                                      �?                                              "@                                       @                                                      @                                      @      �?                                       @      �?                                              �?                                       @                                              @                                                      �?      <@      &@      �?                              2@      &@      �?                              .@      @                                      .@      �?                                      $@                                              @      �?                                      @                                              �?      �?                                              �?                                      �?                                                      @                                      @      @      �?                                      @                                      @              �?                              @                                                              �?                      �?      $@                                      �?      @                                               @                                      �?      �?                                              �?                                      �?                                                      @                              &@      @      0@                              $@              �?                              @                                              @              �?                                              �?                              @                                              �?      @      .@                              �?      @       @                              �?       @       @                              �?      �?                                      �?                                                      �?                                              �?       @                                      �?      @                                              @                                      �?                                                      @                                       @                                                      @                              �?      @                                              @                                      �?                                              @      0@      ,@      (@      2@      @      �?      *@      *@      @      &@       @      �?      *@      $@      @      &@       @              @      @       @      &@       @              @      @       @      @       @              @      �?               @       @              @                       @       @              @                      �?      �?                                      �?      �?                                      �?                                                      �?              @                                                                      �?      �?                                              �?                                      �?                              �?                                               @       @      �?                                       @      �?                                              �?                                       @                                       @                                                               @              �?      "@      @      �?                      �?      @      @      �?                              @                                      �?      �?      @      �?                      �?              @      �?                      �?              �?      �?                      �?                                                              �?      �?                                              �?                                      �?                                              @                                      �?                                              @       @                                      @                                               @       @                                       @                                                       @                                              @      �?                                      �?      �?                                      �?                                                      �?                                       @                               @      @      �?       @      @      @              @      �?       @      @      @                      �?      @      @      @                              @      �?                                      @                                                      �?                              �?      �?      @      @                              �?      @      @                              �?      �?      @                              �?      �?                                              �?                                      �?                                                              @                                       @                              �?              @                              �?                                                              @                      @               @                                               @                              @                                       @                                              @      @      &@      4@      ?@      .@      @      @      &@      4@      (@      @       @      �?       @      3@      @      @      �?              @      @      @       @                      @      @               @                      @      �?               @                      @                                                      �?               @                                               @                              �?                                              @                      �?              �?      @      @              �?              �?      @                                      �?                              �?                      @                      �?                                                                      @                                                      @              �?      �?      �?      (@              �?      �?      �?      �?                              �?              �?                                              �?                              �?                                                      �?                                                              (@              �?                                              �?                              (@                       @       @      @      �?       @       @               @      @      �?      �?       @                       @      �?      �?       @                       @                                                      �?      �?       @                              �?                                                      �?       @                                      �?                                                       @               @      �?                                       @                                                      �?                               @                              @               @                                                                              @                                              3@      $@                                      2@      @                                      2@                                                      @                                      �?      @                                      �?                                                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hKhNhJO�#hG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KK߅�h��B�0         x       &             �?�,����?�            `u@       C                    �?q*�k�?i             e@                           �?��¦��?8            �T@                           �?2Y�Qo��?             ;@                           �?X�<ݚ�?             2@                           @������?	             .@       
                    �?r�q��?             (@       	                    @�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?������������������������       �                     �?                           @�q�q�?             @������������������������       �                     �?������������������������       �                      @              !             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?                            �?|	�%���?             "@              (             �?      �?              @������������������������       �                     �?������������������������       �                     �?                           �?؇���X�?             @������������������������       �                     @                           @�q�q�?             @������������������������       �                      @������������������������       �                     �?       .                    @@��CM?�?%            �K@       #                    @Ǻ����?             9@       "                    �?      �?              @       !                      @r�q��?             @                            �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @$       +                    �?J,�ѳ�?             1@%       (                    �?j�V���?             &@&       '                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @)       *                    �?      �?              @������������������������       �                     @������������������������       �                     �?,       -                    �?�q�q�?             @������������������������       �                      @������������������������       �                     @/       >                    �?�H�7�&�?             >@0       5                    �?(������?             9@1       4                    �?�θ�?             *@2       3       #             �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @6       ;                    @�������?             (@7       :                    �?ףp=
�?             $@8       9                    �?؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @<       =                    @      �?              @������������������������       �                     �?������������������������       �                     �??       @                    �?{�G�z�?             @������������������������       �                      @A       B       	             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @D       U                     �?}�P�z�?1            �U@E       R                    �?����?            �@@F       M                    �?��E���?             ;@G       H                    �?&���^B�?             2@������������������������       �                     $@I       L       (             �?      �?              @J       K                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @N       O                    �?X�<ݚ�?             "@������������������������       �                     @P       Q                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?S       T                    �?�q�q�?             @������������������������       �                     @������������������������       �                      @V       s                    @���y��?"             K@W       p                    �?����R�?            �D@X       o                    @�.k���?             A@Y       n                    @      �?             @@Z       e                    �?���ؓ�?             ?@[       d                    �?�LQ�1	�?             7@\       ]                    @�C��2(�?             6@������������������������       �                     1@^       c                    �?���Q��?             @_       b                    �?      �?             @`       a                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     �?f       m                    �?      �?              @g       h                     @0�����?             @������������������������       �                     �?i       j                    �?r�q��?             @������������������������       �                     @k       l                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @q       r       "             �?؇���X�?             @������������������������       �                     @������������������������       �                     �?t       u       '             �?$�q-�?             *@������������������������       �                     "@v       w                    @      �?             @������������������������       �                     �?������������������������       �                     @y       �                    �?nΪ�>k�?i            �e@z       �                    �?\�O�Mc�?`            �c@{       �       (             �?�	B�~�?            �A@|       �                    �?ĳ���o�?             >@}       �                    �?r
^N���?             <@~       �                    �?0�����?             2@       �                     �?�IєX�?             1@�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �        	             (@������������������������       �                     �?�       �       '             �?      �?             $@������������������������       �                     @�       �       #             �?r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    @_�fѸ��?J            @^@�       �                    �?����z�?#            �O@�       �                     @      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?l�(�|�?!            �N@�       �       
             �?�MbX9�?             I@�       �                    @�eP*L��?             F@�       �       "             �?P���Q�?             D@������������������������       �                     ?@�       �                    �?�<ݚ�?             "@�       �                     �?����X�?             @�       �                    �?r�q��?             @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                    @      �?             @������������������������       �                      @������������������������       �                      @�       �       #             �?�8��8��?             @������������������������       �                      @�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �?�x?r���?             &@�       �                    �?�Q����?             @������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?�q�q�?             @������������������������       �                     @�       �       !             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    @K������?'             M@�       �                    �?c�ee��?            �H@�       �                     @��}��?            �E@�       �                    �?      �?              @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     �?�       �                    @      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?������?            �A@�       �                    �?؇���X�?             @������������������������       �                     @������������������������       �                     �?�       �                    �? �Cc}�?             <@������������������������       �                     1@�       �                    �?���!pc�?	             &@������������������������       �                     @�       �                    �?      �?             @������������������������       �                      @�       �       !             �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?r�q��?             @������������������������       �                     �?������������������������       �                     @�       �       !             �?��E���?             "@�       �                    @����X�?             @������������������������       �                      @������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �       )             �?�M�]��?	             1@�       �                    �?      �?             (@�       �                    �?�����H�?             "@������������������������       �                      @������������������������       �                     �?�       �                     @�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    @���Q��?             @������������������������       �                     @������������������������       �                      @�t�bh�h)h,K ��h.��R�(KK�KK��h�B�)       �@@      T@      V@     @P@     �H@      ;@      @      @     �C@      I@      G@      8@              �?      6@      2@     �@@       @              �?       @      *@      @      �?                       @      (@      @                                      &@      @                                      $@       @                                      $@      �?                                      $@                                                      �?                                              �?                                      �?       @                                      �?                                                       @                               @      �?                                       @                                                      �?                              �?      @      �?              �?              �?              �?                              �?                                                              �?                                      @                      �?                      @                                               @                      �?                       @                                                                      �?                      ,@      @      =@      @                      "@      @       @      @                      @      �?                                      @      �?                                       @      �?                                       @                                                      �?                                      @                                               @                                               @      @       @      @                       @      �?       @                               @              �?                                              �?                               @                                                      �?      @                                              @                                      �?                                               @              @                               @                                                              @                      @      �?      5@      @                      @      �?      4@      �?                      @              $@                              @               @                                               @                              @                                                               @                                      �?      $@      �?                              �?      "@                                      �?      @                                      �?                                                      @                                              @                                              �?      �?                                      �?                                                      �?                       @              �?       @                                               @                       @              �?                                              �?                               @                              @      @      1@      @@      *@      0@      �?      @      .@      @      @      @      �?      @      .@      @      �?                      @      *@              �?                              $@                                      @      @              �?                              @              �?                                              �?                              @                                      @                                      �?               @      @                                              @                      �?               @                                               @                              �?                                                                               @      @                                              @                                       @              @      �?       @      :@      $@      (@      @      �?       @      :@      "@              @      �?       @      9@      @              �?      �?       @      9@      @              �?      �?      �?      9@      @                                      4@      @                                      4@       @                                      1@                                              @       @                                      @      �?                                      �?      �?                                      �?                                                      �?                                       @                                                      �?                                              �?              �?      �?      �?      @                              �?      �?      @                              �?                                                      �?      @                                              @                                      �?       @                                      �?                                                       @                      �?                                                              �?                               @                                                                      �?      @                                              @                                      �?                                                      �?      (@                                              "@                                      �?      @                                      �?                                                      @      =@     �R@     �H@      .@      @      @      =@     @Q@     �C@      *@      @      @      5@      @      @      �?              �?      5@       @      @      �?              �?      5@      �?      @      �?                      0@      �?              �?                      0@      �?                                      @      �?                                              �?                                      @                                              (@                                                                      �?                      @              @                              @                                              �?              @                                              @                              �?                                                      �?                              �?                                              �?              �?                                              @                                       @      O@      A@      (@      @       @      @      G@      @      @       @              �?              �?                              �?                                                              �?                              @      G@      @      @       @              @     �D@      @               @               @      C@       @               @               @      C@                                              ?@                                       @      @                                       @      @                                      �?      @                                      �?       @                                               @                                      �?                                                      @                                      �?                                                       @                                                       @               @                               @                                                               @              �?      @       @                                               @                              �?      @                                      �?                                                      @                                      �?      @       @      @                      �?      �?              @                                              @                      �?      �?                                      �?                                                      �?                                              @       @                                      @                                              �?       @                                               @                                      �?                                      @      0@      ;@      "@      �?       @      @      0@      9@      @              �?      @      &@      9@      @                       @      @              �?                              @                                       @                      �?                      �?                                              �?                      �?                      �?                                                                      �?                      �?      @      9@      @                      �?      @                                              @                                      �?                                                              9@      @                                      1@                                               @      @                                      @                                              �?      @                                               @                                      �?      �?                                      �?                                                      �?                              @                              �?                                              �?              @                                                       @      @      �?      �?                       @      @                                       @                                                      @                                                      �?      �?                                      �?                                                      �?              @      $@       @                               @       @       @                                       @      �?                                       @                                                      �?                               @              �?                               @                                                              �?                              @       @                                      @                                                       @                        �t�bubhhubh)��}�(hhhhhNhKhKhG        hKhNhJ��^hG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKh��BH4         �       &             �?��7M��?�            `u@       c                    �?&�9A���?y            �f@       "                    �?��0�Q��?`            �a@                           �?9��8���?             B@              "             �?��k����?             :@                           �?8�Z$���?
             *@                            @      �?              @                           @�Q����?             @	       
                     �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @                           @�T�6|��?
             *@                           �?�C��2(�?             &@������������������������       �                      @                             @�q�q�?             @������������������������       �                     �?������������������������       �                      @              
             �?      �?              @������������������������       �                     �?������������������������       �                     �?       !                    �?��Q��?             $@              "             �?      �?              @                           �?z�G�z�?             @������������������������       �                     @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?                            �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @#       :                    @b����{�?E            @Z@$       9                    @\���	�?             C@%       *                    @+�{72Y�?             ;@&       '                    �?�����H�?             "@������������������������       �                     @(       )                      @      �?              @������������������������       �                     �?������������������������       �                     �?+       .                    �?���[���?             2@,       -                    �?      �?             @������������������������       �                      @������������������������       �                      @/       8                    �?X�Cc�?
             ,@0       7                    �?�eP*L��?             &@1       2                    @�q�q�?             "@������������������������       �                     �?3       6                     @      �?              @4       5                    �?؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     &@;       \                    �?����?+            �P@<       S                    �?��<��)�?$            �J@=       P       	             �?N�mL�?            �E@>       O       $             �?�xRvQ��?            �C@?       N                    �?P���� �?             7@@       E       !             �?j�V���?             6@A       D                    @�C��2(�?             &@B       C                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@F       K                    �?Y�����?             &@G       J                    @�q�q�?             @H       I       '             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?L       M                    @      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     0@Q       R       "             �?      �?             @������������������������       �                     @������������������������       �                     �?T       [                    @���(\��?	             $@U       Z                    �?�$I�$I�?             @V       Y                    �?      �?             @W       X                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @]       b                    �?      �?             ,@^       _                    @�<ݚ�?             "@������������������������       �                     �?`       a       
             �?      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     @d       �                    �?�G�z��?             D@e       �                    �?�5?,R�?             B@f       q                    @8,�̂�?             ?@g       p                     @.k��\�?
             1@h       i                    �?     ��?	             0@������������������������       �                      @j       o       #             �?@4և���?             ,@k       l                    @z�G�z�?             @������������������������       �                      @m       n                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     "@������������������������       �                     �?r       y                    �?$I�$I��?	             ,@s       x                    �?      �?             @t       u       )             �?z�G�z�?             @������������������������       �                     @v       w                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?z                           �?      �?              @{       ~                    �?�Q����?             @|       }                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    �?=�c����?h             d@�       �                    �?M��>�?Z             a@�       �                     �?H���I}�?1            @T@�       �                    �?؇���X�?             ,@������������������������       �                     "@�       �                    @���Q��?             @������������������������       �                      @������������������������       �                     @�       �                    �?d� ���?*            �P@�       �                    �?��w?I|�?$            �M@�       �                    �?+�����?             I@�       �                    �?r٣����?            �@@�       �                    �?      �?             @@������������������������       �                     @�       �                    �?؇���X�?             <@�       �                    �?`2U0*��?             9@������������������������       �                     0@�       �                     @�����H�?             "@�       �                     �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     �?�       �                    @:���I�?             1@�       �                    �?�m۶m��?             ,@������������������������       �                      @�       �                    �?�8��8��?             @�       �                    �?      �?             @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                     �?�2�tk~�?             "@�       �       #             �?      �?             @������������������������       �                      @������������������������       �                      @�       �                    �?�Q����?             @�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �       )             �?      �?              @�       �                    @VUUUUU�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �       !             �?��;�9�?)            �K@�       �       $             �?>
ףp=�?             D@�       �                    @c�=��?             ?@�       �                    �?b'vb'v�?             :@�       �                     @�8��8��?             @�       �       )             �?      �?             @������������������������       �                     @������������������������       �                     �?�       �       )             �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?p=
ףp�?             4@�       �                    �?������?             @�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    @.y0��k�?             *@�       �                     �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    @      �?              @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �?h/�����?             "@�       �                    �?����X�?             @������������������������       �                     �?�       �                    @r�q��?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                     @VUUUUU�?             .@�       �                    �?���Q��?             @������������������������       �                     @������������������������       �                      @�       �                    �?p=
ףp�?             $@�       �                    �?�<ݚ�?             "@������������������������       �                     @������������������������       �                      @������������������������       �                     �?�       �                    @n���?             9@�       �                    @�n_Y�K�?             *@�       �                    @      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     "@�       �                    �?      �?             (@������������������������       �                      @�       �                    @ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@�t�bh�h)h,K ��h.��R�(KK�KK��h�B�,        @@     @P@      R@     �U@     �M@      ;@               @     �@@      M@     �L@      9@              @      2@      E@      L@      4@              @      @      2@      $@      �?                       @      ,@      "@      �?                      �?      @       @                              �?      @      @                              �?      �?      @                              �?      �?                                              �?                                      �?                                                              @                                      @                                                      @                              �?      $@      �?      �?                      �?      $@                                               @                                      �?       @                                      �?                                                       @                                                      �?      �?                                              �?                                      �?                      @      �?      @      �?                      @      �?       @      �?                      @      �?                                      @                                              �?      �?                                              �?                                      �?                                                               @      �?                                              �?                                       @                                               @                              �?      .@      8@      G@      3@              �?      .@      4@       @                      �?      .@      "@       @                      �?       @                                              @                                      �?      �?                                      �?                                                      �?                                              @      "@       @                               @               @                               @                                                               @                              @      "@                                      @      @                                      @      @                                      �?                                               @      @                                      �?      @                                              @                                      �?                                              �?                                               @                                                      @                                              &@                                              @      F@      3@                              @     �B@      (@                              @     �@@      @                              @      @@      @                              @      0@      @                               @      0@      @                              �?      $@                                      �?      �?                                              �?                                      �?                                                      "@                                      �?      @      @                              �?       @                                      �?      �?                                      �?                                                      �?                                              �?                                              @      @                                      @                                                      @                              �?                                                      0@                                              �?      @                                              @                                      �?                                      �?      @      @                              �?      @       @                              �?      �?       @                              �?               @                                               @                              �?                                                      �?                                              @                                                      @                                      @      @                                      @       @                                              �?                                      @      �?                                      @                                                      �?                                              @              @      .@      0@      �?      @              @      .@      (@      �?      @              @      .@       @      �?      @              @      *@      �?                              @      *@                                       @                                              �?      *@                                      �?      @                                               @                                      �?       @                                      �?                                                       @                                              "@                                                      �?                                       @      @      �?      @                      �?      �?              @                      �?                      @                                              @                      �?                      �?                      �?                                                                      �?                              �?                                      �?      @      �?                              �?      @      �?                              �?      @                                              @                                      �?                                                              �?                                      @                                              @              �?                              @                                                              �?                              @                      @@     �L@     �C@      =@       @       @      >@     �K@      ;@      4@       @       @      1@      D@      .@      @       @      �?              (@       @                                      "@                                              @       @                                               @                                      @                                      1@      <@      *@      @       @      �?      &@      ;@      (@      @       @      �?      "@      ;@      &@      @                       @      9@                                       @      8@                                      @                                              @      8@                                      �?      8@                                              0@                                      �?       @                                      �?       @                                      �?                                                       @                                              @                                      @                                                      �?                                      �?       @      &@      @                      �?       @      &@                                               @                              �?       @      @                              �?       @      �?                                       @      �?                                              �?                                       @                                      �?                                                               @                                                      @                       @              �?      @       @      �?       @                               @               @                                                                               @                              �?      @              �?                      �?      @                                              @                                      �?                                                                      �?      @      �?      �?                              �?      �?      �?                              �?      �?                                              �?                                      �?                                                              �?                              @                                              *@      .@      (@      ,@              �?      $@      .@       @      @                      @      .@      @      @                      @      .@      @                              @      �?       @                              @              �?                              @                                                              �?                                      �?      �?                                      �?                                                      �?                               @      ,@      @                              �?      @      @                              �?      @                                              @                                      �?                                                              @                              �?      &@      �?                              �?      @                                              @                                      �?                                                      @      �?                                       @      �?                                       @                                                      �?                                      @                                                              @                      @               @       @                      @               @                                              �?                              @              �?                              �?              �?                                              �?                              �?                                              @                                                                       @                      @              @      @              �?      @               @                              @                                                               @                                               @      @              �?                       @      @                                              @                                       @                                                                      �?       @       @      (@      "@                       @       @      "@                               @       @                                               @                                       @                                                              "@                                              @      "@                                       @                                              �?      "@                                      �?                                                      "@                �t�bub�S      hhubh)��}�(hhhhhNhKhKhG        hKhNhJ�	�^hG        hNhG        heK*hfKhgh)h,K ��h.��R�(KK��h�C0              �?       @      @      @      @�t�bhsh�hnC       ���R�h�Kh�h�K*h)h,K ��h.��R�(KK��hn�C       �t�bK��R�}�(hKh�K�h�h)h,K ��h.��R�(KKɅ�h��B�+         t       &             �?���q��?�            `u@       A                    @(�EY� �?h            �d@       0                    �?z3�Vf`�?6            �T@       +                    @��$���?'            �O@       (       "             �?؛bv�X�?!            �J@       !       !             �?}��7�?             F@                           �?)O���?             B@              )             �?_�g����?             6@	                           �?b���i��?	             &@
                           �?      �?              @������������������������       �                     @                           �?      �?             @������������������������       �                      @                             @      �?              @������������������������       �                     �?������������������������       �                     �?                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @                           �?j�V���?             &@                           �?�<ݚ�?             "@������������������������       �                     @                             @�q�q�?             @������������������������       �                     �?������������������������       �                      @                           @      �?              @������������������������       �                     �?������������������������       �                     �?                           �?؇���X�?             ,@������������������������       �                     $@                            @      �?             @������������������������       �                      @������������������������       �                      @"       '                    �?      �?              @#       &                    �?�q�q�?             @$       %                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                      @)       *                    @�<ݚ�?             "@������������������������       �                     @������������������������       �                      @,       -       
             �?p=
ףp�?             $@������������������������       �                      @.       /                    �?      �?              @������������������������       �                     @������������������������       �                     �?1       >                    �?���.�?             3@2       9                    �?����2�?             .@3       8       '             �?      �?              @4       7       $             �?�8��8��?             @5       6                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @:       =                    @0�����?             @;       <                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @?       @                    �?      �?             @������������������������       �                     �?������������������������       �                     @B       [                    �?���Z�_�?2            �T@C       R                    @��|�5��?            �G@D       M                    �?�[")�i�?
             7@E       H                     @������?             *@F       G                    �?և���X�?             @������������������������       �                     @������������������������       �                     @I       L                    @      �?             @J       K                     �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @N       Q                    �?z�G�z�?             $@O       P       )             �?�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @S       X                    @      �?             8@T       W                     @���N8�?             5@U       V                    @ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?������������������������       �                     &@Y       Z                    @�q�q�?             @������������������������       �                     �?������������������������       �                      @\       e                    @�Kh/��?             B@]       ^                    @�������?             8@������������������������       �                     @_       d                    @:/����?             5@`       a                    �?�KM�]�?             3@������������������������       �        	             0@b       c                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @f       g                    �?�q�q�?	             (@������������������������       �                     �?h       i                    �?�eP*L��?             &@������������������������       �                     �?j       k                    �?      �?             $@������������������������       �                     �?l       s                    @X�<ݚ�?             "@m       n       !             �?�q�q�?             @������������������������       �                     �?o       r                    �?���Q��?             @p       q                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @u       �                    @�ۦ�qA�?e             f@v       {                    �?�}n&P��?1            �V@w       z                    �?AA�?             5@x       y                    �?�}�+r��?             3@������������������������       �        
             2@������������������������       �                     �?������������������������       �                      @|       �       $             �?�:�����?%            @Q@}       �                    @�ƣ�]:�?            �I@~       �                    �?��0{9�?            �G@       �                    �?�}�+r��?             C@�       �       
             �?�?�|�?            �B@������������������������       �                     9@�       �       )             �?�8��8��?             (@������������������������       �                     @�       �                    @      �?              @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                    �?X�<ݚ�?             "@�       �                     �?      �?              @�       �                    �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                    @      �?             @������������������������       �                      @������������������������       �                      @�       �                    �?n�����?
             2@�       �                    �?������?             @�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �?Y�����?             &@�       �                    �?      �?             @������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �?��1"���?4            �U@�       �       $             �?b�H�U��?#             M@�       �                    �?��7���?            �G@������������������������       �                     �?�       �                    �?B�>�)
�?             G@�       �                    @�r����?             >@������������������������       �                     .@�       �                    �?������?	             .@������������������������       �                     @�       �                    @X�<ݚ�?             "@�       �                    �?����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @�       �                    �?     ��?             0@�       �                    @z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    @���!pc�?             &@������������������������       �                      @������������������������       �                     @�       �                    @�C��2(�?             &@�       �                    �?�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                    �?���Q��?             @������������������������       �                      @������������������������       �                     @�       �                    �?����5�?             =@�       �                    �?�q�q�?             (@������������������������       �                      @�       �                    �?�z�G��?             $@������������������������       �                     @�       �       "             �?���Q��?             @������������������������       �                      @������������������������       �                     @�       �       
             �?ҳ�wY;�?
             1@������������������������       �                      @�       �                     @�q�q�?             "@������������������������       �                     @������������������������       �                     @�t�bh�h)h,K ��h.��R�(KK�KK��h�B�%       �E@     �P@     �V@     �Q@      K@      1@      @      @      B@     �H@     �J@      .@              @      <@      5@      7@      @              �?      ;@      1@      .@      @              �?      ;@      .@       @       @              �?      ;@       @      @       @              �?      7@      @      @       @              �?      &@      @      @       @              �?      @      @      @                      �?       @      @      �?                                      @                              �?       @              �?                               @                                      �?                      �?                      �?                                                                      �?                              �?               @                              �?                                                               @                               @              �?       @                      @                       @                      @                                              �?                       @                      �?                                                                       @                      �?              �?                              �?                                                              �?                              (@               @                              $@                                               @               @                               @                                                               @                              @      @                                       @      @                                      �?      @                                      �?                                                      @                                      �?                                               @                                                      @       @                                      @                                                       @                                       @      @      �?                               @                                                      @      �?                                      @                                                      �?               @      �?      @       @      @              �?      �?      @       @      �?                              @      @      �?                               @      @      �?                               @              �?                               @                                                              �?                                      @                                       @                              �?      �?              @                      �?      �?                                      �?                                                      �?                                                              @                      �?                              @              �?                                                                              @      @      @       @      <@      >@       @      @      @      @      &@      5@      @      @      @      @      &@                      @      @      @      @                      @      @                                      @                                                      @                                                      @      @                                      @      �?                                      @                                                      �?                                               @                       @                       @                       @                      @                       @                                                                      @                                              @                                                      5@      @                                      4@      �?                                      "@      �?                                      "@                                                      �?                                      &@                                              �?       @                                      �?                                                       @                      @      1@      "@      @                      @      1@       @                              @                                               @      1@       @                               @      1@                                              0@                                       @      �?                                       @                                                      �?                                                       @                                              @      @                                      �?                                              @      @                                      �?                                              @      @                                      �?                                              @      @                                      @       @                                      �?                                              @       @                                      @      �?                                              �?                                      @                                                      �?                                              @     �B@     �N@     �K@      5@      �?       @      ?@      G@      @      @               @      2@      �?                               @      2@      �?                                      2@                                                      �?                                                                               @      *@     �F@      @      @                      @      D@       @       @                      @      D@                                       @      B@                                      �?      B@                                              9@                                      �?      &@                                              @                                      �?      @                                      �?      �?                                      �?                                                      �?                                              @                                      �?                                              @      @                                      @      @                                       @      @                                              @                                       @                                              @                                                      �?                                                       @       @                                       @                                                       @                      @      @      @      @                              �?      @      @                              �?      @                                      �?                                                      @                                                      @                      @      @      �?                              �?      @      �?                                      @                                      �?              �?                              �?                                                              �?                              @                                              @      .@     �H@      0@      �?              �?       @      C@      $@      �?              �?      @      A@      @      �?                                              �?              �?      @      A@      @                                      :@      @                                      .@                                              &@      @                                      @                                              @      @                                      @       @                                               @                                      @                                                       @                      �?      @       @      @                      �?      @                                              @                                      �?                                                               @      @                                       @                                                      @                              @      @      @                              @       @                                      @                                                       @                                               @      @                                       @                                                      @                      @      @      &@      @                      @      @                                       @                                              @      @                                              @                                      @       @                                               @                                      @                                                              &@      @                                       @                                              @      @                                              @                                      @                        �t�bubhhubehhub.